
module Connect4 ( CLK, NRST, start, G, O, LED_PIN, C4_OUT );
  input [3:0] G;
  input [3:0] O;
  output [23:0] LED_PIN;
  output [1:0] C4_OUT;
  input CLK, NRST, start;
  wire   N683, N684, N689, N690, N692, N693, N694, N695, N696, N698, N699,
         N700, N701, N702, N704, N705, N706, N707, N708, N716, N717, N718,
         N719, N720, N722, N723, N724, N725, N726, N740, N741, N742, N743,
         N744, N837, N838, N839, N840, N842, N843, N844, N845, N846, N850,
         N851, N852, N855, N856, N857, N858, N860, N861, N862, N863, N864,
         N873, N874, N875, N876, N940, N941, N942, N952, N953, N954, N956,
         N957, N958, N959, N960, N964, N965, N966, N968, N969, N970, N971,
         N972, N975, N976, N977, N978, N980, N981, N982, N983, N984, N987,
         N988, N989, N990, N993, N994, N995, N996, N998, N999, N1000, N1001,
         N1002, N1004, N1005, N1006, N1007, N1008, N1010, N1011, N1012, N1013,
         N1014, N1016, N1017, N1018, N1019, N1020, N1022, N1023, N1024, N1025,
         N1026, N1029, N1030, N1031, N1032, N1034, N1035, N1036, N1037, N1038,
         N1040, N1041, N1042, N1043, N1044, N1046, N1047, N1048, N1049, N1050,
         N1053, N1054, N1055, N1056, N1059, N1060, N1061, N1062, N1066, N1067,
         N1068, N1072, N1073, N1074, N1077, N1078, N1079, N1080, N1082, N1083,
         N1084, N1085, N1086, N1107, N1108, N1109, N1110, N1112, N1113, N1114,
         N1115, N1116, N1120, N1121, N1122, N1125, N1126, N1127, N1128, N1130,
         N1131, N1132, N1133, N1134, N1138, N1139, N1140, N1143, N1144, N1145,
         N1146, N1148, N1149, N1150, N1151, N1152, N1156, N1157, N1158, N1161,
         N1162, N1163, N1164, N1167, N1168, N1169, N1170, N1172, N1173, N1174,
         N1175, N1176, N1180, N1181, N1182, N1184, N1185, N1186, N1187, N1188,
         N1191, N1192, N1193, N1194, N1197, N1198, N1199, N1200, N1203, N1204,
         N1205, N1206, N1207, N1208, N1210, N1211, N1212, N1215, N1216, N1217,
         N1218, N1220, N1221, N1222, N1223, N1224, N1228, N1229, N1230, N1233,
         N1234, N1235, N1236, N1240, N1241, N1242, N1244, N1245, N1246, N1247,
         N1248, N1252, N1253, N1254, N1256, N1257, N1258, N1259, N1260, N1263,
         N1264, N1265, N1266, \Col_Fill[7][31] , \Col_Fill[7][30] ,
         \Col_Fill[7][29] , \Col_Fill[7][28] , \Col_Fill[7][27] ,
         \Col_Fill[7][26] , \Col_Fill[7][25] , \Col_Fill[7][24] ,
         \Col_Fill[7][23] , \Col_Fill[7][22] , \Col_Fill[7][21] ,
         \Col_Fill[7][20] , \Col_Fill[7][19] , \Col_Fill[7][18] ,
         \Col_Fill[7][17] , \Col_Fill[7][16] , \Col_Fill[7][15] ,
         \Col_Fill[7][14] , \Col_Fill[7][13] , \Col_Fill[7][12] ,
         \Col_Fill[7][11] , \Col_Fill[7][10] , \Col_Fill[7][9] ,
         \Col_Fill[7][8] , \Col_Fill[7][7] , \Col_Fill[7][6] ,
         \Col_Fill[7][5] , \Col_Fill[7][4] , \Col_Fill[7][3] ,
         \Col_Fill[7][2] , \Col_Fill[7][1] , \Col_Fill[7][0] ,
         \Col_Fill[6][31] , \Col_Fill[6][30] , \Col_Fill[6][29] ,
         \Col_Fill[6][28] , \Col_Fill[6][27] , \Col_Fill[6][26] ,
         \Col_Fill[6][25] , \Col_Fill[6][24] , \Col_Fill[6][23] ,
         \Col_Fill[6][22] , \Col_Fill[6][21] , \Col_Fill[6][20] ,
         \Col_Fill[6][19] , \Col_Fill[6][18] , \Col_Fill[6][17] ,
         \Col_Fill[6][16] , \Col_Fill[6][15] , \Col_Fill[6][14] ,
         \Col_Fill[6][13] , \Col_Fill[6][12] , \Col_Fill[6][11] ,
         \Col_Fill[6][10] , \Col_Fill[6][9] , \Col_Fill[6][8] ,
         \Col_Fill[6][7] , \Col_Fill[6][6] , \Col_Fill[6][5] ,
         \Col_Fill[6][4] , \Col_Fill[6][3] , \Col_Fill[6][2] ,
         \Col_Fill[6][1] , \Col_Fill[6][0] , \Col_Fill[5][31] ,
         \Col_Fill[5][30] , \Col_Fill[5][29] , \Col_Fill[5][28] ,
         \Col_Fill[5][27] , \Col_Fill[5][26] , \Col_Fill[5][25] ,
         \Col_Fill[5][24] , \Col_Fill[5][23] , \Col_Fill[5][22] ,
         \Col_Fill[5][21] , \Col_Fill[5][20] , \Col_Fill[5][19] ,
         \Col_Fill[5][18] , \Col_Fill[5][17] , \Col_Fill[5][16] ,
         \Col_Fill[5][15] , \Col_Fill[5][14] , \Col_Fill[5][13] ,
         \Col_Fill[5][12] , \Col_Fill[5][11] , \Col_Fill[5][10] ,
         \Col_Fill[5][9] , \Col_Fill[5][8] , \Col_Fill[5][7] ,
         \Col_Fill[5][6] , \Col_Fill[5][5] , \Col_Fill[5][4] ,
         \Col_Fill[5][3] , \Col_Fill[5][2] , \Col_Fill[5][1] ,
         \Col_Fill[5][0] , \Col_Fill[4][31] , \Col_Fill[4][30] ,
         \Col_Fill[4][29] , \Col_Fill[4][28] , \Col_Fill[4][27] ,
         \Col_Fill[4][26] , \Col_Fill[4][25] , \Col_Fill[4][24] ,
         \Col_Fill[4][23] , \Col_Fill[4][22] , \Col_Fill[4][21] ,
         \Col_Fill[4][20] , \Col_Fill[4][19] , \Col_Fill[4][18] ,
         \Col_Fill[4][17] , \Col_Fill[4][16] , \Col_Fill[4][15] ,
         \Col_Fill[4][14] , \Col_Fill[4][13] , \Col_Fill[4][12] ,
         \Col_Fill[4][11] , \Col_Fill[4][10] , \Col_Fill[4][9] ,
         \Col_Fill[4][8] , \Col_Fill[4][7] , \Col_Fill[4][6] ,
         \Col_Fill[4][5] , \Col_Fill[4][4] , \Col_Fill[4][3] ,
         \Col_Fill[4][2] , \Col_Fill[4][1] , \Col_Fill[4][0] ,
         \Col_Fill[3][31] , \Col_Fill[3][30] , \Col_Fill[3][29] ,
         \Col_Fill[3][28] , \Col_Fill[3][27] , \Col_Fill[3][26] ,
         \Col_Fill[3][25] , \Col_Fill[3][24] , \Col_Fill[3][23] ,
         \Col_Fill[3][22] , \Col_Fill[3][21] , \Col_Fill[3][20] ,
         \Col_Fill[3][19] , \Col_Fill[3][18] , \Col_Fill[3][17] ,
         \Col_Fill[3][16] , \Col_Fill[3][15] , \Col_Fill[3][14] ,
         \Col_Fill[3][13] , \Col_Fill[3][12] , \Col_Fill[3][11] ,
         \Col_Fill[3][10] , \Col_Fill[3][9] , \Col_Fill[3][8] ,
         \Col_Fill[3][7] , \Col_Fill[3][6] , \Col_Fill[3][5] ,
         \Col_Fill[3][4] , \Col_Fill[3][3] , \Col_Fill[3][2] ,
         \Col_Fill[3][1] , \Col_Fill[3][0] , \Col_Fill[2][31] ,
         \Col_Fill[2][30] , \Col_Fill[2][29] , \Col_Fill[2][28] ,
         \Col_Fill[2][27] , \Col_Fill[2][26] , \Col_Fill[2][25] ,
         \Col_Fill[2][24] , \Col_Fill[2][23] , \Col_Fill[2][22] ,
         \Col_Fill[2][21] , \Col_Fill[2][20] , \Col_Fill[2][19] ,
         \Col_Fill[2][18] , \Col_Fill[2][17] , \Col_Fill[2][16] ,
         \Col_Fill[2][15] , \Col_Fill[2][14] , \Col_Fill[2][13] ,
         \Col_Fill[2][12] , \Col_Fill[2][11] , \Col_Fill[2][10] ,
         \Col_Fill[2][9] , \Col_Fill[2][8] , \Col_Fill[2][7] ,
         \Col_Fill[2][6] , \Col_Fill[2][5] , \Col_Fill[2][4] ,
         \Col_Fill[2][3] , \Col_Fill[2][2] , \Col_Fill[2][1] ,
         \Col_Fill[2][0] , \Col_Fill[1][31] , \Col_Fill[1][30] ,
         \Col_Fill[1][29] , \Col_Fill[1][28] , \Col_Fill[1][27] ,
         \Col_Fill[1][26] , \Col_Fill[1][25] , \Col_Fill[1][24] ,
         \Col_Fill[1][23] , \Col_Fill[1][22] , \Col_Fill[1][21] ,
         \Col_Fill[1][20] , \Col_Fill[1][19] , \Col_Fill[1][18] ,
         \Col_Fill[1][17] , \Col_Fill[1][16] , \Col_Fill[1][15] ,
         \Col_Fill[1][14] , \Col_Fill[1][13] , \Col_Fill[1][12] ,
         \Col_Fill[1][11] , \Col_Fill[1][10] , \Col_Fill[1][9] ,
         \Col_Fill[1][8] , \Col_Fill[1][7] , \Col_Fill[1][6] ,
         \Col_Fill[1][5] , \Col_Fill[1][4] , \Col_Fill[1][3] ,
         \Col_Fill[1][2] , \Col_Fill[1][1] , \Col_Fill[1][0] ,
         \Col_Fill[0][31] , \Col_Fill[0][30] , \Col_Fill[0][29] ,
         \Col_Fill[0][28] , \Col_Fill[0][27] , \Col_Fill[0][26] ,
         \Col_Fill[0][25] , \Col_Fill[0][24] , \Col_Fill[0][23] ,
         \Col_Fill[0][22] , \Col_Fill[0][21] , \Col_Fill[0][20] ,
         \Col_Fill[0][19] , \Col_Fill[0][18] , \Col_Fill[0][17] ,
         \Col_Fill[0][16] , \Col_Fill[0][15] , \Col_Fill[0][14] ,
         \Col_Fill[0][13] , \Col_Fill[0][12] , \Col_Fill[0][11] ,
         \Col_Fill[0][10] , \Col_Fill[0][9] , \Col_Fill[0][8] ,
         \Col_Fill[0][7] , \Col_Fill[0][6] , \Col_Fill[0][5] ,
         \Col_Fill[0][4] , \Col_Fill[0][3] , \Col_Fill[0][2] ,
         \Col_Fill[0][1] , \Col_Fill[0][0] , \GFill[63][0] , \GFill[62][0] ,
         \GFill[61][0] , \GFill[60][0] , \GFill[59][0] , \GFill[58][0] ,
         \GFill[57][0] , \GFill[56][0] , \GFill[55][0] , \GFill[54][0] ,
         \GFill[53][0] , \GFill[52][0] , \GFill[51][0] , \GFill[50][0] ,
         \GFill[49][0] , \GFill[48][0] , \GFill[47][0] , \GFill[46][0] ,
         \GFill[45][0] , \GFill[44][0] , \GFill[43][0] , \GFill[42][0] ,
         \GFill[41][0] , \GFill[40][0] , \GFill[39][0] , \GFill[38][0] ,
         \GFill[37][0] , \GFill[36][0] , \GFill[35][0] , \GFill[34][0] ,
         \GFill[33][0] , \GFill[32][0] , \GFill[31][0] , \GFill[30][0] ,
         \GFill[29][0] , \GFill[28][0] , \GFill[27][0] , \GFill[26][0] ,
         \GFill[25][0] , \GFill[24][0] , \GFill[23][0] , \GFill[22][0] ,
         \GFill[21][0] , \GFill[20][0] , \GFill[19][0] , \GFill[18][0] ,
         \GFill[17][0] , \GFill[16][0] , \GFill[15][0] , \GFill[14][0] ,
         \GFill[13][0] , \GFill[12][0] , \GFill[11][0] , \GFill[10][0] ,
         \GFill[9][0] , \GFill[8][0] , \GFill[7][0] , \GFill[6][0] ,
         \GFill[5][0] , \GFill[4][0] , \GFill[3][0] , \GFill[2][0] ,
         \GFill[1][0] , \GFill[0][0] , \OFill[63][0] , \OFill[62][0] ,
         \OFill[61][0] , \OFill[60][0] , \OFill[59][0] , \OFill[58][0] ,
         \OFill[57][0] , \OFill[56][0] , \OFill[55][0] , \OFill[54][0] ,
         \OFill[53][0] , \OFill[52][0] , \OFill[51][0] , \OFill[50][0] ,
         \OFill[49][0] , \OFill[48][0] , \OFill[47][0] , \OFill[46][0] ,
         \OFill[45][0] , \OFill[44][0] , \OFill[43][0] , \OFill[42][0] ,
         \OFill[41][0] , \OFill[40][0] , \OFill[39][0] , \OFill[38][0] ,
         \OFill[37][0] , \OFill[36][0] , \OFill[35][0] , \OFill[34][0] ,
         \OFill[33][0] , \OFill[32][0] , \OFill[31][0] , \OFill[30][0] ,
         \OFill[29][0] , \OFill[28][0] , \OFill[27][0] , \OFill[26][0] ,
         \OFill[25][0] , \OFill[24][0] , \OFill[23][0] , \OFill[22][0] ,
         \OFill[21][0] , \OFill[20][0] , \OFill[19][0] , \OFill[18][0] ,
         \OFill[17][0] , \OFill[16][0] , \OFill[15][0] , \OFill[14][0] ,
         \OFill[13][0] , \OFill[12][0] , \OFill[11][0] , \OFill[10][0] ,
         \OFill[9][0] , \OFill[8][0] , \OFill[7][0] , \OFill[6][0] ,
         \OFill[5][0] , \OFill[4][0] , \OFill[3][0] , \OFill[2][0] ,
         \OFill[1][0] , \OFill[0][0] , N1293, N1294, N1295, N1300, N1301,
         N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311,
         N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321,
         N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331,
         N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341,
         N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351,
         N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361,
         N1362, N1367, N1368, N1371, N1404, N1405, N1406, N1407, N1408, N1409,
         N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, N1419,
         N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, N1429,
         N1430, N1431, N1432, N1433, N1434, N1435, N1439, N1440, N1441, N1442,
         N1443, N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452,
         N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462,
         N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1472, N1473,
         N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483,
         N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493,
         N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503,
         N1506, N1507, N1508, N1509, N1510, N1515, N1516, N1517, N1518, N1519,
         N1520, N1521, N1522, N1523, N1524, N1526, N1527, N1528, N1529, N1530,
         N1560, N1836, N1837, N1838, N1843, N1844, N1845, N1846, N1847, N1848,
         N1849, N1850, N1851, N1852, N1853, N1854, N1855, N1856, N1857, N1858,
         N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868,
         N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878,
         N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1886, N1887, N1888,
         N1889, N1890, N1891, N1892, N1893, N1894, N1895, N1896, N1897, N1898,
         N1899, N1900, N1901, N1902, N1903, N1904, N1905, N1910, N1911, N1914,
         N1947, N1948, N1949, N1950, N1951, N1952, N1953, N1954, N1955, N1956,
         N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1964, N1965, N1966,
         N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976,
         N1977, N1978, N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989,
         N1990, N1991, N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999,
         N2000, N2001, N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009,
         N2010, N2011, N2012, N2013, N2015, N2016, N2017, N2018, N2019, N2020,
         N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030,
         N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040,
         N2041, N2042, N2043, N2044, N2045, N2046, N2049, N2050, N2051, N2052,
         N2053, N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066,
         N2067, N2070, N2071, N2072, N2073, N2103, N2629, N2630, N2631, N2632,
         N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642,
         N2643, N2644, N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652,
         N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662,
         N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672,
         N2673, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2713, N2714,
         N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2723, N2724,
         N2725, N2726, N2727, N2728, N2729, N2730, N2731, N2732, N2733, N2734,
         N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744,
         N2745, N2746, N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754,
         N2755, N2756, N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764,
         N2765, N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774,
         N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784,
         N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794,
         N2795, N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804,
         N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814,
         N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824,
         N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834,
         N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844,
         N2845, N2846, N2847, N2848, N2849, N3008, N3040, N3194, N3195, N3196,
         N3200, N3285, N3317, N3349, N3351, N3472, N3504, N3505, N3599, N3631,
         N3758, N3760, N3988, N4020, N4021, N4092, N4124, N4156, N4229, N4261,
         N4293, N4294, N4295, N4297, N4368, N4400, N4432, N4434, N4436, N4571,
         N4572, N4573, N4602, N4603, N4708, N4709, N4728, N4781, N4813, N4845,
         N4847, N4849, N4855, N4920, N4952, N4984, N4985, N4986, N4988, N5058,
         N5090, N5122, N5124, N5246, N5278, N5310, N5400, N5432, N5464, N5555,
         N5587, N5619, N5710, N5742, N5774, N5837, N5869, N5901, N5964, N5996,
         N6028, N6226, N6258, N6290, N6362, N6394, N6426, N6499, N6531, N6563,
         N6638, N6670, N6702, N6777, N6809, N6841, N6914, N6946, N6978, N7051,
         N7083, N7115, N7190, N7222, N7254, N7328, N7360, N7392, n1654, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1696, n1703, n1708, n1709, n1718, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1761, n1762, n1803,
         n1804, n1805, n1846, n1847, n1848, n1890, n1931, n1932, n1973, n1974,
         n1975, n2016, n2017, n2018, n2060, n2102, n2103, n2145, n2146, n2230,
         n2231, n2244, n2273, n2274, n2315, n2316, n2358, n2399, n2400, n2413,
         n2414, n2443, n2444, n2486, n2487, n2528, n2529, n2570, n2571, n2612,
         n2613, n2654, n2655, n2696, n2697, n2738, n2739, n2780, n2781, n2794,
         n2824, n2825, n2910, n2911, n2952, n2953, n2994, n2995, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3121, n3122, n3163, n3164, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3321,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n25099, n25100, n25101, n25102, n25103,
         n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
         n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n26379, n26380, n26381, n26382, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26392, n26393, n26394, n26395, n26396, n26397, n26398, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27659, n27660, n27661, n27662, n27663,
         n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671,
         n27672, n27673, n27674, n27675, n27676, n27677, n27678, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28939, n28940, n28941, n28942, n28943,
         n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
         n28952, n28953, n28954, n28955, n28956, n28957, n28958, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n30219, n30220, n30221, n30222, n30223,
         n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231,
         n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30859,
         n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
         n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
         n30876, n30877, n30878, n31499, n31500, n31501, n31502, n31503,
         n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511,
         n31512, n31513, n31514, n31515, n31516, n31517, n31518, n32139,
         n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
         n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
         n32156, n32157, n32158, n32779, n32780, n32781, n32782, n32783,
         n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791,
         n32792, n32793, n32794, n32795, n32796, n32797, n32798, n33419,
         n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
         n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435,
         n33436, n33437, n33438, n34059, n34060, n34061, n34062, n34063,
         n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071,
         n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34699,
         n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707,
         n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715,
         n34716, n34717, n34718, n35339, n35340, n35341, n35342, n35343,
         n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351,
         n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35979,
         n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987,
         n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
         n35996, n35997, n35998, n36619, n36620, n36621, n36622, n36623,
         n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631,
         n36632, n36633, n36634, n36635, n36636, n36637, n36638, n37259,
         n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267,
         n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275,
         n37276, n37277, n37278, n37899, n37900, n37901, n37902, n37903,
         n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911,
         n37912, n37913, n37914, n37915, n37916, n37917, n37918, n38539,
         n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547,
         n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555,
         n38556, n38557, n38558, n39179, n39180, n39181, n39182, n39183,
         n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191,
         n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39819,
         n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827,
         n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
         n39836, n39837, n39838, n40459, n40460, n40461, n40462, n40463,
         n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471,
         n40472, n40473, n40474, n40475, n40476, n40477, n40478, n41099,
         n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107,
         n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115,
         n41116, n41117, n41118, n41739, n41740, n41741, n41742, n41743,
         n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751,
         n41752, n41753, n41754, n41755, n41756, n41757, n41758, n42379,
         n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387,
         n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395,
         n42396, n42397, n42398, n43019, n43020, n43021, n43022, n43023,
         n43024, n43025, n43026, n43027, n43028, n43029, n43030, n43031,
         n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43659,
         n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
         n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675,
         n43676, n43677, n43678, n44299, n44300, n44301, n44302, n44303,
         n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311,
         n44312, n44313, n44314, n44315, n44316, n44317, n44318, n44939,
         n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
         n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955,
         n44956, n44957, n44958, n45579, n45580, n45581, n45582, n45583,
         n45584, n45585, n45586, n45587, n45588, n45589, n45590, n45591,
         n45592, n45593, n45594, n45595, n45596, n45597, n45598, n48139,
         n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147,
         n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155,
         n48156, n48157, n48158, n48779, n48780, n48781, n48782, n48783,
         n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791,
         n48792, n48793, n48794, n48795, n48796, n48797, n48798, n49419,
         n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427,
         n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435,
         n49436, n49437, n49438, n50059, n50060, n50061, n50062, n50063,
         n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071,
         n50072, n50073, n50074, n50075, n50076, n50077, n50078, n50699,
         n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707,
         n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715,
         n50716, n50717, n50718, n51339, n51340, n51341, n51342, n51343,
         n51344, n51345, n51346, n51347, n51348, n51349, n51350, n51351,
         n51352, n51353, n51354, n51355, n51356, n51357, n51358, n51979,
         n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987,
         n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995,
         n51996, n51997, n51998, n52619, n52620, n52621, n52622, n52623,
         n52624, n52625, n52626, n52627, n52628, n52629, n52630, n52631,
         n52632, n52633, n52634, n52635, n52636, n52637, n52638, n53259,
         n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267,
         n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275,
         n53276, n53277, n53278, n53899, n53900, n53901, n53902, n53903,
         n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911,
         n53912, n53913, n53914, n53915, n53916, n53917, n53918, n54539,
         n54540, n54541, n54542, n54543, n54544, n54545, n54546, n54547,
         n54548, n54549, n54550, n54551, n54552, n54553, n54554, n54555,
         n54556, n54557, n54558, n55179, n55180, n55181, n55182, n55183,
         n55184, n55185, n55186, n55187, n55188, n55189, n55190, n55191,
         n55192, n55193, n55194, n55195, n55196, n55197, n55198, n55819,
         n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827,
         n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835,
         n55836, n55837, n55838, n56459, n56460, n56461, n56462, n56463,
         n56464, n56465, n56466, n56467, n56468, n56469, n56470, n56471,
         n56472, n56473, n56474, n56475, n56476, n56477, n56478, n57099,
         n57100, n57101, n57102, n57103, n57104, n57105, n57106, n57107,
         n57108, n57109, n57110, n57111, n57112, n57113, n57114, n57115,
         n57116, n57117, n57118, n57739, n57740, n57741, n57742, n57743,
         n57744, n57745, n57746, n57747, n57748, n57749, n57750, n57751,
         n57752, n57753, n57754, n57755, n57756, n57757, n57758, n58379,
         n58380, n58381, n58382, n58383, n58384, n58385, n58386, n58387,
         n58388, n58389, n58390, n58391, n58392, n58393, n58394, n58395,
         n58396, n58397, n58398, n59019, n59020, n59021, n59022, n59023,
         n59024, n59025, n59026, n59027, n59028, n59029, n59030, n59031,
         n59032, n59033, n59034, n59035, n59036, n59037, n59038, n59659,
         n59660, n59661, n59662, n59663, n59664, n59665, n59666, n59667,
         n59668, n59669, n59670, n59671, n59672, n59673, n59674, n59675,
         n59676, n59677, n59678, n60299, n60300, n60301, n60302, n60303,
         n60304, n60305, n60306, n60307, n60308, n60309, n60310, n60311,
         n60312, n60313, n60314, n60315, n60316, n60317, n60318, n60939,
         n60940, n60941, n60942, n60943, n60944, n60945, n60946, n60947,
         n60948, n60949, n60950, n60951, n60952, n60953, n60954, n60955,
         n60956, n60957, n60958, n61579, n61580, n61581, n61582, n61583,
         n61584, n61585, n61586, n61587, n61588, n61589, n61590, n61591,
         n61592, n61593, n61594, n61595, n61596, n61597, n61598, n62219,
         n62220, n62221, n62222, n62223, n62224, n62225, n62226, n62227,
         n62228, n62229, n62230, n62231, n62232, n62233, n62234, n62235,
         n62236, n62237, n62238, n62859, n62860, n62861, n62862, n62863,
         n62864, n62865, n62866, n62867, n62868, n62869, n62870, n62871,
         n62872, n62873, n62874, n62875, n62876, n62877, n62878, n63499,
         n63500, n63501, n63502, n63503, n63504, n63505, n63506, n63507,
         n63508, n63509, n63510, n63511, n63512, n63513, n63514, n63515,
         n63516, n63517, n63518, n64139, n64140, n64141, n64142, n64143,
         n64144, n64145, n64146, n64147, n64148, n64149, n64150, n64151,
         n64152, n64153, n64154, n64155, n64156, n64157, n64158, n64779,
         n64780, n64781, n64782, n64783, n64784, n64785, n64786, n64787,
         n64788, n64789, n64790, n64791, n64792, n64793, n64794, n64795,
         n64796, n64797, n64798, \sub_143_2_cf/carry[2] ,
         \sub_143_2_cf/carry[3] , \sub_143_2_cf/carry[4] ,
         \sub_143_2_cf/carry[5] , \sub_143_2_cf/carry[6] , N11532, N11531,
         N11530, N7278, N7277, N11526, N11525, N11524, N7266, N11544, N11543,
         N11542, N5008, N5007, N11538, N11537, N11536, N4996, N4858, N4857,
         N11514, N11513, N11512, N7152, N7151, N11508, N11507, N11506, N7140,
         N4882, N4881, N11520, N11519, N11518, N4870, N4731, N4730, N11496,
         N11495, N11494, N4719, N4718, N11490, N11489, N11488, N7013, N4743,
         N4606, N4605, N11472, N11471, N11470, N4594, N4593, N11466, N11465,
         N11464, N4582, N4581, N11460, N11459, N11458, N4469, N4468, N11436,
         N11435, N11434, N4457, N4456, N11430, N11429, N11428, N4445, N4444,
         N4330, N4329, N11412, N11411, N11410, N4318, N4317, N6576, N11394,
         N11393, N11392, N4306, N11406, N11405, N11404, N4191, N4190, N6449,
         N6448, N11376, N11375, N11374, N6437, N11370, N11369, N11368, N4179,
         N4178, N11388, N11387, N11386, N4167, N11382, N11381, N11380, N11346,
         N11345, N11344, N6312, N6311, N11340, N11339, N11338, N6300, N11334,
         N11333, N11332, N11363, N11362, N4042, N4041, N11357, N11356, N4030,
         N11351, N11350, N3900, N3899, N11322, N11321, N11320, N3638, N3637,
         N11292, N11291, N11290, N11286, N11285, N11284, N3511, N3510, N11268,
         N11267, N11266, N11262, N11261, N11260, N11256, N11255, N11254, N3402,
         N3401, N3400, N3396, N3395, N3384, N3383, N3382, N3378, N3377, N3366,
         N3365, N3364, N3360, N3359, N3229, N3228, N3227, N3223, N3222, N3211,
         N3210, N3209, N3205, N3204, N5517, N5516, N5515, N5511, N3247, N3246,
         N3245, N3241, N11206, N11205, N11204, N11203, N11202, N11216, N11215,
         N11214, N11213, N11212, N3056, N3055, N3054, N3050, N3049, N5362,
         N5361, N5360, N5356, N5355, N5344, N5343, N5342, N5338, N3092, N3091,
         N3090, N3086, N3085, N3074, N3073, N3072, N3068, N1403, N1380, N1379,
         N1378, N1377, N1376, N1946, N1923, N1922, N1921, N1920, N1919, n807,
         N5208, N5207, N5206, N5190, N5189, N5188, N5184, N5183, N5172, N5171,
         N5170, N5166, N2938, N2937, N2936, N2920, N2919, N2914, N2913, N2902,
         N2901, N2896, \add_1_root_add_157_3/carry[2] , \r11555/carry[5] ,
         \r11554/carry[5] , \r11553/carry[5] , \r12189/carry[3] ,
         \r12189/carry[4] , \r12189/carry[5] , \r12187/carry[5] ,
         \r13449/carry[5] , \r13448/carry[5] ,
         \add_1_root_add_0_root_sub_325_4_cf/carry[5] ,
         \add_1_root_add_0_root_sub_325_8_cf/carry[5] ,
         \add_1_root_add_0_root_sub_325_12_cf/carry[5] ,
         \add_1_root_add_0_root_sub_397_8_cf/carry[3] ,
         \add_1_root_add_0_root_sub_397_8_cf/carry[4] ,
         \add_1_root_add_0_root_sub_328_4_cf/carry[4] ,
         \add_1_root_add_0_root_sub_328_8_cf/carry[2] ,
         \add_1_root_add_0_root_sub_328_8_cf/carry[5] ,
         \add_1_root_add_0_root_sub_400_4_cf/carry[5] ,
         \add_1_root_add_0_root_sub_400_8_cf/carry[5] ,
         \add_1_root_add_0_root_sub_331_4_cf/carry[4] ,
         \add_1_root_add_0_root_sub_403_4_cf/carry[5] , \add_342_5/carry[5] ,
         \add_414_5/carry[5] , \add_345_3/carry[5] , \add_345_5/carry[5] ,
         \add_417_3/carry[5] , \add_417_5/carry[5] , \add_348/carry[5] ,
         \add_348_3/carry[5] , \add_420/carry[5] , \add_420_3/carry[5] ,
         \add_1_root_add_126_3/carry[2] , \r2195/n5 , \r2195/n4 , \r2195/n3 ,
         \r2182/n5 , \r2182/n4 , \r2182/n3 , \sub_171_2_cf/carry[2] ,
         \sub_171_2_cf/carry[3] , \sub_171_2_cf/carry[4] ,
         \sub_171_2_cf/carry[5] , \sub_171_2_cf/carry[6] ,
         \sub_171_2_cf/carry[7] , \sub_171_2_cf/carry[8] ,
         \sub_171_2_cf/carry[9] , \sub_171_2_cf/carry[10] , \r30598/carry[3] ,
         \r30598/carry[4] , \r30598/carry[5] , \r31195/carry[5] ,
         \r33598/carry[4] , \r33598/carry[5] , \r35376/carry[5] ,
         \r35965/carry[5] , \r39563/carry[5] , \r40165/carry[5] ,
         \r41369/carry[4] , \sub_1_root_sub_0_root_sub_167_2/A[4] ,
         \sub_1_root_sub_0_root_sub_136_2/A[4] , n65419, n65420, n65421,
         n65422, n65423, n65424, n65425, n65426, n65427, n65428, n65429,
         n65430, n65431, n65432, n65433, n65434, n65435, n65436, n65437,
         n65438, n65439, n65440, n65441, n65442, n65443, n65444, n65445,
         n65446, n65447, n65448, n65449, n65450, n65451, n65452, n65453,
         n65454, n65455, n65456, n65457, n65458, n65459, n65460, n65461,
         n65462, n65463, n65464, n65465, n65466, n65467, n65468, n65469,
         n65470, n65471, n65472, n65473, n65474, n65475, n65476, n65477,
         n65478, n65479, n65480, n65481, n65482, n65483, n65484, n65485,
         n65486, n65487, n65488, n65489, n65490, n65491, n65492, n65493,
         n65494, n65495, n65496, n65497, n65498, n65499, n65500, n65501,
         n65502, n65503, n65504, n65505, n65506, n65507, n65508, n65509,
         n65510, n65511, n65512, n65513, n65514, n65515, n65516, n65517,
         n65518, n65519, n65520, n65521, n65522, n65523, n65524, n65525,
         n65526, n65527, n65528, n65529, n65530, n65531, n65532, n65533,
         n65534, n65535, n65536, n65537, n65538, n65539, n65540, n65541,
         n65542, n65543, n65544, n65545, n65546, n65547, n65548, n65549,
         n65550, n65551, n65552, n65553, n65554, n65555, n65556, n65557,
         n65558, n65559, n65560, n65561, n65562, n65563, n65564, n65565,
         n65566, n65567, n65568, n65569, n65570, n65571, n65572, n65573,
         n65574, n65575, n65576, n65577, n65578, n65579, n65580, n65581,
         n65582, n65583, n65584, n65585, n65586, n65587, n65588, n65589,
         n65590, n65591, n65592, n65593, n65594, n65595, n65596, n65597,
         n65598, n65599, n65600, n65601, n65602, n65603, n65604, n65605,
         n65606, n65607, n65608, n65609, n65610, n65611, n65612, n65613,
         n65614, n65615, n65616, n65617, n65618, n65619, n65620, n65621,
         n65622, n65623, n65624, n65625, n65626, n65627, n65628, n65629,
         n65630, n65631, n65632, n65633, n65634, n65635, n65636, n65637,
         n65638, n65639, n65640, n65641, n65642, n65643, n65644, n65645,
         n65646, n65647, n65648, n65649, n65650, n65651, n65652, n65653,
         n65654, n65655, n65656, n65657, n65658, n65659, n65660, n65661,
         n65662, n65663, n65664, n65665, n65666, n65667, n65668, n65669,
         n65670, n65671, n65672, n65673, n65674, n65675, n65676, n65677,
         n65678, n65679, n65680, n65681, n65682, n65683, n65684, n65685,
         n65686, n65687, n65688, n65689, n65690, n65691, n65692, n65693,
         n65694, n65695, n65696, n65697, n65698, n65699, n65700, n65701,
         n65702, n65703, n65704, n65705, n65706, n65707, n65708, n65709,
         n65710, n65711, n65712, n65713, n65714, n65715, n65716, n65717,
         n65718, n65719, n65720, n65721, n65722, n65723, n65724, n65725,
         n65726, n65727, n65728, n65729, n65730, n65731, n65732, n65733,
         n65734, n65735, n65736, n65737, n65738, n65739, n65740, n65741,
         n65742, n65743, n65744, n65745, n65746, n65747, n65748, n65749,
         n65750, n65751, n65752, n65753, n65754, n65755, n65756, n65757,
         n65758, n65759, n65760, n65761, n65762, n65763, n65764, n65765,
         n65766, n65767, n65768, n65769, n65770, n65771, n65772, n65773,
         n65774, n65775, n65776, n65777, n65778, n65779, n65780, n65781,
         n65782, n65783, n65784, n65785, n65786, n65787, n65788, n65789,
         n65790, n65791, n65792, n65793, n65794, n65795, n65796, n65797,
         n65798, n65799, n65800, n65801, n65802, n65803, n65804, n65805,
         n65806, n65807, n65808, n65809, n65810, n65811, n65812, n65813,
         n65814, n65815, n65816, n65817, n65818, n65819, n65820, n65821,
         n65822, n65823, n65824, n65825, n65826, n65827, n65828, n65829,
         n65830, n65831, n65832, n65833, n65834, n65835, n65836, n65837,
         n65838, n65839, n65840, n65841, n65842, n65843, n65844, n65845,
         n65846, n65847, n65848, n65849, n65850, n65851, n65852, n65853,
         n65854, n65855, n65856, n65857, n65858, n65859, n65860, n65861,
         n65862, n65863, n65864, n65865, n65866, n65867, n65868, n65869,
         n65870, n65871, n65872, n65873, n65874, n65875, n65876, n65877,
         n65878, n65879, n65880, n65881, n65882, n65883, n65884, n65885,
         n65886, n65887, n65888, n65889, n65890, n65891, n65892, n65893,
         n65894, n65895, n65896, n65897, n65898, n65899, n65900, n65901,
         n65902, n65903, n65904, n65905, n65906, n65907, n65908, n65909,
         n65910, n65911, n65912, n65913, n65914, n65915, n65916, n65917,
         n65918, n65919, n65920, n65921, n65922, n65923, n65924, n65925,
         n65926, n65927, n65928, n65929, n65930, n65931, n65932, n65933,
         n65934, n65935, n65936, n65937, n65938, n65939, n65940, n65941,
         n65942, n65943, n65944, n65945, n65946, n65947, n65948, n65949,
         n65950, n65951, n65952, n65953, n65954, n65955, n65956, n65957,
         n65958, n65959, n65960, n65961, n65962, n65963, n65964, n65965,
         n65966, n65967, n65968, n65969, n65970, n65971, n65972, n65973,
         n65974, n65975, n65976, n65977, n65978, n65979, n65980, n65981,
         n65982, n65983, n65984, n65985, n65986, n65987, n65988, n65989,
         n65990, n65991, n65992, n65993, n65994, n65995, n65996, n65997,
         n65998, n65999, n66000, n66001, n66002, n66003, n66004, n66005,
         n66006, n66007, n66008, n66009, n66010, n66011, n66012, n66013,
         n66014, n66015, n66016, n66017, n66018, n66019, n66020, n66021,
         n66022, n66023, n66024, n66025, n66026, n66027, n66028, n66029,
         n66030, n66031, n66032, n66033, n66034, n66035, n66036, n66037,
         n66038, n66039, n66040, n66041, n66042, n66043, n66044, n66045,
         n66046, n66047, n66048, n66049, n66050, n66051, n66052, n66053,
         n66054, n66055, n66056, n66057, n66058, n66059, n66060, n66061,
         n66062, n66063, n66064, n66065, n66066, n66067, n66068, n66069,
         n66070, n66071, n66072, n66073, n66074, n66075, n66076, n66077,
         n66078, n66079, n66080, n66081, n66082, n66083, n66084, n66085,
         n66086, n66087, n66088, n66089, n66090, n66091, n66092, n66093,
         n66094, n66095, n66096, n66097, n66098, n66099, n66100, n66101,
         n66102, n66103, n66104, n66105, n66106, n66107, n66108, n66109,
         n66110, n66111, n66112, n66113, n66114, n66115, n66116, n66117,
         n66118, n66119, n66120, n66121, n66122, n66123, n66124, n66125,
         n66126, n66127, n66128, n66129, n66130, n66131, n66132, n66133,
         n66134, n66135, n66136, n66137, n66138, n66139, n66140, n66141,
         n66142, n66143, n66144, n66145, n66146, n66147, n66148, n66149,
         n66150, n66151, n66152, n66153, n66154, n66155, n66156, n66157,
         n66158, n66159, n66160, n66161, n66162, n66163, n66164, n66165,
         n66166, n66167, n66168, n66169, n66170, n66171, n66172, n66173,
         n66174, n66175, n66176, n66177, n66178, n66179, n66180, n66181,
         n66182, n66183, n66184, n66185, n66186, n66187, n66188, n66189,
         n66190, n66191, n66192, n66193, n66194, n66195, n66196, n66197,
         n66198, n66199, n66200, n66201, n66202, n66203, n66204, n66205,
         n66206, n66207, n66208, n66209, n66210, n66211, n66212, n66213,
         n66214, n66215, n66216, n66217, n66218, n66219, n66220, n66221,
         n66222, n66223, n66224, n66225, n66226, n66227, n66228, n66229,
         n66230, n66231, n66232, n66233, n66234, n66235, n66236, n66237,
         n66238, n66239, n66240, n66241, n66242, n66243, n66244, n66245,
         n66246, n66247, n66248, n66249, n66250, n66251, n66252, n66253,
         n66254, n66255, n66256, n66257, n66258, n66259, n66260, n66261,
         n66262, n66263, n66264, n66265, n66266, n66267, n66268, n66269,
         n66270, n66271, n66272, n66273, n66274, n66275, n66276, n66277,
         n66278, n66279, n66280, n66281, n66282, n66283, n66284, n66285,
         n66286, n66287, n66288, n66289, n66290, n66291, n66292, n66293,
         n66294, n66295, n66296, n66297, n66298, n66299, n66300, n66301,
         n66302, n66303, n66304, n66305, n66306, n66307, n66308, n66309,
         n66310, n66311, n66312, n66313, n66314, n66315, n66316, n66317,
         n66318, n66319, n66320, n66321, n66322, n66323, n66324, n66325,
         n66326, n66327, n66328, n66329, n66330, n66331, n66332, n66333,
         n66334, n66335, n66336, n66337, n66338, n66339, n66340, n66341,
         n66342, n66343, n66344, n66345, n66346, n66347, n66348, n66349,
         n66350, n66351, n66352, n66353, n66354, n66355, n66356, n66357,
         n66358, n66359, n66360, n66361, n66362, n66363, n66364, n66365,
         n66366, n66367, n66368, n66369, n66370, n66371, n66372, n66373,
         n66374, n66375, n66376, n66377, n66378, n66379, n66380, n66381,
         n66382, n66383, n66384, n66385, n66386, n66387, n66388, n66389,
         n66390, n66391, n66392, n66393, n66394, n66395, n66396, n66397,
         n66398, n66399, n66400, n66401, n66402, n66403, n66404, n66405,
         n66406, n66407, n66408, n66409, n66410, n66411, n66412, n66413,
         n66414, n66415, n66416, n66417, n66418, n66419, n66420, n66421,
         n66422, n66423, n66424, n66425, n66426, n66427, n66428, n66429,
         n66430, n66431, n66432, n66433, n66434, n66435, n66436, n66437,
         n66438, n66439, n66440, n66441, n66442, n66443, n66444, n66445,
         n66446, n66447, n66448, n66449, n66450, n66451, n66452, n66453,
         n66454, n66455, n66456, n66457, n66458, n66459, n66460, n66461,
         n66462, n66463, n66464, n66465, n66466, n66467, n66468, n66469,
         n66470, n66471, n66472, n66473, n66474, n66475, n66476, n66477,
         n66478, n66479, n66480, n66481, n66482, n66483, n66484, n66485,
         n66486, n66487, n66488, n66489, n66490, n66491, n66492, n66493,
         n66494, n66495, n66496, n66497, n66498, n66499, n66500, n66501,
         n66502, n66503, n66504, n66505, n66506, n66507, n66508, n66509,
         n66510, n66511, n66512, n66513, n66514, n66515, n66516, n66517,
         n66518, n66519, n66520, n66521, n66522, n66523, n66524, n66525,
         n66526, n66527, n66528, n66529, n66530, n66531, n66532, n66533,
         n66534, n66535, n66536, n66537, n66538, n66539, n66540, n66541,
         n66542, n66543, n66544, n66545, n66546, n66547, n66548, n66549,
         n66550, n66551, n66552, n66553, n66554, n66555, n66556, n66557,
         n66558, n66559, n66560, n66561, n66562, n66563, n66564, n66565,
         n66566, n66567, n66568, n66569, n66570, n66571, n66572, n66573,
         n66574, n66575, n66576, n66577, n66578, n66579, n66580, n66581,
         n66582, n66583, n66584, n66585, n66586, n66587, n66588, n66589,
         n66590, n66591, n66592, n66593, n66594, n66595, n66596, n66597,
         n66598, n66599, n66600, n66601, n66602, n66603, n66604, n66605,
         n66606, n66607, n66608, n66609, n66610, n66611, n66612, n66613,
         n66614, n66615, n66616, n66617, n66618, n66619, n66620, n66621,
         n66622, n66623, n66624, n66625, n66626, n66627, n66628, n66629,
         n66630, n66631, n66632, n66633, n66634, n66635, n66636, n66637,
         n66638, n66639, n66640, n66641, n66642, n66643, n66644, n66645,
         n66646, n66647, n66648, n66649, n66650, n66651, n66652, n66653,
         n66654, n66655, n66656, n66657, n66658, n66659, n66660, n66661,
         n66662, n66663, n66664, n66665, n66666, n66667, n66668, n66669,
         n66670, n66671, n66672, n66673, n66674, n66675, n66676, n66677,
         n66678, n66679, n66680, n66681, n66682, n66683, n66684, n66685,
         n66686, n66687, n66688, n66689, n66690, n66691, n66692, n66693,
         n66694, n66695, n66696, n66697, n66698, n66699, n66700, n66701,
         n66702, n66703, n66704, n66705, n66706, n66707, n66708, n66709,
         n66710, n66711, n66712, n66713, n66714, n66715, n66716, n66717,
         n66718, n66719, n66720, n66721, n66722, n66723, n66724, n66725,
         n66726, n66727, n66728, n66729, n66730, n66731, n66732, n66733,
         n66734, n66735, n66736, n66737, n66738, n66739, n66740, n66741,
         n66742, n66743, n66744, n66745, n66746, n66747, n66748, n66749,
         n66750, n66751, n66752, n66753, n66754, n66755, n66756, n66757,
         n66758, n66759, n66760, n66761, n66762, n66763, n66764, n66765,
         n66766, n66767, n66768, n66769, n66770, n66771, n66772, n66773,
         n66774, n66775, n66776, n66777, n66778, n66779, n66780, n66781,
         n66782, n66783, n66784, n66785, n66786, n66787, n66788, n66789,
         n66790, n66791, n66792, n66793, n66794, n66795, n66796, n66797,
         n66798, n66799, n66800, n66801, n66802, n66803, n66804, n66805,
         n66806, n66807, n66808, n66809, n66810, n66811, n66812, n66813,
         n66814, n66815, n66816, n66817, n66818, n66819, n66820, n66821,
         n66822, n66823, n66824, n66825, n66826, n66827, n66828, n66829,
         n66830, n66831, n66832, n66833, n66834, n66835, n66836, n66837,
         n66838, n66839, n66840, n66841, n66842, n66843, n66844, n66845,
         n66846, n66847, n66848, n66849, n66850, n66851, n66852, n66853,
         n66854, n66855, n66856, n66857, n66858, n66859, n66860, n66861,
         n66862, n66863, n66864, n66865, n66866, n66867, n66868, n66869,
         n66870, n66871, n66872, n66873, n66874, n66875, n66876, n66877,
         n66878, n66879, n66880, n66881, n66882, n66883, n66884;
  wire   [1:0] state;
  wire   [1:0] next_state;
  wire   [3:0] G_play;
  wire   [3:0] O_play;
  wire   [31:0] m;
  wire   [31:0] n;
  wire   [10:1] \sub_174_2_cf/carry ;
  wire   [31:2] \add_168/carry ;
  wire   [32:0] \sub_157_S2_2/carry ;
  wire   [31:2] \add_137/carry ;
  wire   [32:0] \sub_126_S2_2/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_297_3/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_297_6/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_297_9/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_369_3/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_369_6/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_369_9/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_300_5/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_300_8/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_372_5/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_372_8/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_303_7/carry ;
  wire   [5:1] \add_0_root_sub_0_root_sub_375_7/carry ;
  wire   [5:1] \r11558/carry ;
  wire   [5:1] \r11557/carry ;
  wire   [5:1] \r11556/carry ;
  wire   [5:1] \r12191/carry ;
  wire   [5:1] \r12190/carry ;
  wire   [5:1] \r12188/carry ;
  wire   [5:2] \r13451/carry ;
  wire   [5:1] \r13450/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_325_4_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_325_8_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_325_12_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_397_4_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_397_8_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_397_12_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_328_4_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_328_8_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_400_4_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_400_8_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_331_4_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_403_4_cf/carry ;
  wire   [5:2] \sub_345_9_cf/carry ;
  wire   [5:2] \sub_417_9_cf/carry ;
  wire   [5:2] \sub_348_6_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_348_9_cf/carry ;
  wire   [5:1] \add_1_root_add_0_root_sub_348_9_cf/carry ;
  wire   [5:2] \sub_420_6_cf/carry ;
  wire   [5:1] \add_0_root_add_0_root_sub_420_9_cf/carry ;
  wire   [10:0] \sub_171_b0/carry ;
  wire   [5:1] \r30599/carry ;
  wire   [5:2] \r31196/carry ;
  wire   [5:1] \r31798/carry ;
  wire   [5:1] \r32400/carry ;
  wire   [5:2] \r32997/carry ;
  wire   [5:1] \r32996/carry ;
  wire   [5:1] \r33599/carry ;
  wire   [10:1] \sub_140_2_cf/carry ;
  wire   [10:0] \sub_140_b0/carry ;
  wire   [5:1] \r34787/carry ;
  wire   [5:1] \r34786/carry ;
  wire   [5:1] \r36567/carry ;
  wire   [5:1] \r37169/carry ;
  wire   [5:1] \r37771/carry ;
  wire   [5:1] \r38360/carry ;
  wire   [5:1] \r38962/carry ;
  wire   [5:1] \r39564/carry ;
  wire   [5:1] \r40166/carry ;
  wire   [5:1] \r40768/carry ;
  wire   [5:1] \r41370/carry ;

  XNR22 U6167 ( .A(N1837), .B(n3177), .Q(N690) );
  XNR22 U6170 ( .A(N1294), .B(n3178), .Q(N684) );
  OAI222 U6215 ( .A(n65533), .B(n3217), .C(n65522), .D(n3218), .Q(N2849) );
  OAI212 U6216 ( .A(n66394), .B(n65590), .C(n65569), .Q(N2848) );
  OAI212 U6218 ( .A(n3219), .B(n3220), .C(n65569), .Q(N2847) );
  OAI212 U6219 ( .A(n3220), .B(n3221), .C(n65569), .Q(N2846) );
  OAI212 U6220 ( .A(n3220), .B(n3222), .C(n65569), .Q(N2845) );
  OAI212 U6221 ( .A(n3220), .B(n3223), .C(n66568), .Q(N2844) );
  OAI212 U6222 ( .A(n3220), .B(n3224), .C(n65569), .Q(N2843) );
  OAI212 U6223 ( .A(n3220), .B(n3225), .C(n66568), .Q(N2842) );
  OAI212 U6224 ( .A(n3220), .B(n3226), .C(n66568), .Q(N2841) );
  OAI212 U6225 ( .A(n3220), .B(n3227), .C(n66568), .Q(N2840) );
  OAI212 U6227 ( .A(n3219), .B(n3228), .C(n66568), .Q(N2839) );
  OAI212 U6228 ( .A(n3221), .B(n3228), .C(n66568), .Q(N2838) );
  OAI212 U6229 ( .A(n3222), .B(n3228), .C(n66568), .Q(N2837) );
  OAI212 U6230 ( .A(n3223), .B(n3228), .C(n65568), .Q(N2836) );
  OAI212 U6231 ( .A(n3224), .B(n3228), .C(n65567), .Q(N2835) );
  OAI212 U6232 ( .A(n3225), .B(n3228), .C(n65567), .Q(N2834) );
  OAI212 U6233 ( .A(n3226), .B(n3228), .C(n66568), .Q(N2833) );
  OAI212 U6234 ( .A(n3227), .B(n3228), .C(n66568), .Q(N2832) );
  OAI212 U6236 ( .A(n3219), .B(n3229), .C(n65568), .Q(N2831) );
  OAI212 U6237 ( .A(n3221), .B(n3229), .C(n65567), .Q(N2830) );
  OAI212 U6238 ( .A(n3222), .B(n3229), .C(n65568), .Q(N2829) );
  OAI212 U6239 ( .A(n3223), .B(n3229), .C(n66568), .Q(N2828) );
  OAI212 U6240 ( .A(n3224), .B(n3229), .C(n66568), .Q(N2827) );
  OAI212 U6241 ( .A(n3225), .B(n3229), .C(n65568), .Q(N2826) );
  OAI212 U6242 ( .A(n3226), .B(n3229), .C(n65567), .Q(N2825) );
  OAI212 U6243 ( .A(n3227), .B(n3229), .C(n65567), .Q(N2824) );
  OAI212 U6245 ( .A(n3219), .B(n3230), .C(n65568), .Q(N2823) );
  OAI212 U6246 ( .A(n3221), .B(n3230), .C(n65568), .Q(N2822) );
  OAI212 U6247 ( .A(n3222), .B(n3230), .C(n65568), .Q(N2821) );
  OAI212 U6248 ( .A(n3223), .B(n3230), .C(n65568), .Q(N2820) );
  OAI212 U6249 ( .A(n3224), .B(n3230), .C(n65568), .Q(N2819) );
  OAI212 U6250 ( .A(n3225), .B(n3230), .C(n65568), .Q(N2818) );
  OAI212 U6251 ( .A(n3226), .B(n3230), .C(n65568), .Q(N2817) );
  OAI212 U6252 ( .A(n3227), .B(n3230), .C(n65568), .Q(N2816) );
  OAI212 U6254 ( .A(n3219), .B(n3231), .C(n65568), .Q(N2815) );
  OAI212 U6255 ( .A(n3221), .B(n3231), .C(n65568), .Q(N2814) );
  OAI212 U6256 ( .A(n3222), .B(n3231), .C(n65568), .Q(N2813) );
  OAI212 U6257 ( .A(n3223), .B(n3231), .C(n65568), .Q(N2812) );
  OAI212 U6258 ( .A(n3224), .B(n3231), .C(n65568), .Q(N2811) );
  OAI212 U6259 ( .A(n3225), .B(n3231), .C(n65568), .Q(N2810) );
  OAI212 U6260 ( .A(n3226), .B(n3231), .C(n65568), .Q(N2809) );
  OAI212 U6261 ( .A(n3227), .B(n3231), .C(n65568), .Q(N2808) );
  OAI212 U6263 ( .A(n3219), .B(n3232), .C(n65568), .Q(N2807) );
  OAI212 U6264 ( .A(n3221), .B(n3232), .C(n65568), .Q(N2806) );
  OAI212 U6265 ( .A(n3222), .B(n3232), .C(n65568), .Q(N2805) );
  OAI212 U6266 ( .A(n3223), .B(n3232), .C(n65568), .Q(N2804) );
  OAI212 U6267 ( .A(n3224), .B(n3232), .C(n65568), .Q(N2803) );
  OAI212 U6268 ( .A(n3225), .B(n3232), .C(n65567), .Q(N2802) );
  OAI212 U6269 ( .A(n3226), .B(n3232), .C(n65567), .Q(N2801) );
  OAI212 U6270 ( .A(n3227), .B(n3232), .C(n65567), .Q(N2800) );
  OAI212 U6272 ( .A(n3219), .B(n3233), .C(n65567), .Q(N2799) );
  OAI212 U6273 ( .A(n3221), .B(n3233), .C(n65567), .Q(N2798) );
  OAI212 U6274 ( .A(n3222), .B(n3233), .C(n65567), .Q(N2797) );
  OAI212 U6275 ( .A(n3223), .B(n3233), .C(n65567), .Q(N2796) );
  OAI212 U6276 ( .A(n3224), .B(n3233), .C(n65567), .Q(N2795) );
  OAI212 U6277 ( .A(n3225), .B(n3233), .C(n65567), .Q(N2794) );
  OAI212 U6278 ( .A(n3226), .B(n3233), .C(n65567), .Q(N2793) );
  OAI212 U6279 ( .A(n3227), .B(n3233), .C(n65567), .Q(N2792) );
  OAI212 U6281 ( .A(n3219), .B(n3234), .C(n65567), .Q(N2791) );
  OAI212 U6283 ( .A(n3221), .B(n3234), .C(n65567), .Q(N2790) );
  OAI212 U6285 ( .A(n3222), .B(n3234), .C(n65567), .Q(N2789) );
  OAI212 U6287 ( .A(n3223), .B(n3234), .C(n65567), .Q(N2788) );
  OAI212 U6289 ( .A(n3224), .B(n3234), .C(n65567), .Q(N2787) );
  OAI212 U6291 ( .A(n3225), .B(n3234), .C(n65567), .Q(N2786) );
  OAI212 U6293 ( .A(n3226), .B(n3234), .C(n65567), .Q(N2785) );
  OAI212 U6295 ( .A(n3227), .B(n3234), .C(n65567), .Q(N2784) );
  OAI212 U6308 ( .A(n3245), .B(n3246), .C(n65567), .Q(N2783) );
  OAI212 U6309 ( .A(n3246), .B(n3247), .C(n65567), .Q(N2782) );
  OAI212 U6310 ( .A(n3246), .B(n3248), .C(n65568), .Q(N2781) );
  OAI212 U6311 ( .A(n3246), .B(n3249), .C(n65567), .Q(N2780) );
  OAI212 U6312 ( .A(n3246), .B(n3250), .C(n65568), .Q(N2779) );
  OAI212 U6313 ( .A(n3246), .B(n3251), .C(n65567), .Q(N2778) );
  OAI212 U6314 ( .A(n3246), .B(n3252), .C(n65568), .Q(N2777) );
  OAI212 U6315 ( .A(n3246), .B(n3253), .C(n65567), .Q(N2776) );
  OAI212 U6317 ( .A(n3245), .B(n3254), .C(n65568), .Q(N2775) );
  OAI212 U6318 ( .A(n3247), .B(n3254), .C(n65567), .Q(N2774) );
  OAI212 U6319 ( .A(n3248), .B(n3254), .C(n65568), .Q(N2773) );
  OAI212 U6320 ( .A(n3249), .B(n3254), .C(n65567), .Q(N2772) );
  OAI212 U6321 ( .A(n3250), .B(n3254), .C(n65568), .Q(N2771) );
  OAI212 U6322 ( .A(n3251), .B(n3254), .C(n65567), .Q(N2770) );
  OAI212 U6323 ( .A(n3252), .B(n3254), .C(n65568), .Q(N2769) );
  OAI212 U6324 ( .A(n3253), .B(n3254), .C(n65567), .Q(N2768) );
  OAI212 U6326 ( .A(n3245), .B(n3255), .C(n65568), .Q(N2767) );
  OAI212 U6327 ( .A(n3247), .B(n3255), .C(n65567), .Q(N2766) );
  OAI212 U6328 ( .A(n3248), .B(n3255), .C(n65568), .Q(N2765) );
  OAI212 U6329 ( .A(n3249), .B(n3255), .C(n65567), .Q(N2764) );
  OAI212 U6330 ( .A(n3250), .B(n3255), .C(n65568), .Q(N2763) );
  OAI212 U6331 ( .A(n3251), .B(n3255), .C(n65567), .Q(N2762) );
  OAI212 U6332 ( .A(n3252), .B(n3255), .C(n65568), .Q(N2761) );
  OAI212 U6333 ( .A(n3253), .B(n3255), .C(n65568), .Q(N2760) );
  OAI212 U6335 ( .A(n3245), .B(n3256), .C(n65567), .Q(N2759) );
  OAI212 U6336 ( .A(n3247), .B(n3256), .C(n66568), .Q(N2758) );
  OAI212 U6337 ( .A(n3248), .B(n3256), .C(n66568), .Q(N2757) );
  OAI212 U6338 ( .A(n3249), .B(n3256), .C(n65568), .Q(N2756) );
  OAI212 U6339 ( .A(n3250), .B(n3256), .C(n65567), .Q(N2755) );
  OAI212 U6340 ( .A(n3251), .B(n3256), .C(n65568), .Q(N2754) );
  OAI212 U6341 ( .A(n3252), .B(n3256), .C(n65568), .Q(N2753) );
  OAI212 U6342 ( .A(n3253), .B(n3256), .C(n65567), .Q(N2752) );
  OAI212 U6344 ( .A(n3245), .B(n3257), .C(n65567), .Q(N2751) );
  OAI212 U6345 ( .A(n3247), .B(n3257), .C(n65568), .Q(N2750) );
  OAI212 U6346 ( .A(n3248), .B(n3257), .C(n65567), .Q(N2749) );
  OAI212 U6347 ( .A(n3249), .B(n3257), .C(n65568), .Q(N2748) );
  OAI212 U6348 ( .A(n3250), .B(n3257), .C(n65568), .Q(N2747) );
  OAI212 U6349 ( .A(n3251), .B(n3257), .C(n65567), .Q(N2746) );
  OAI212 U6350 ( .A(n3252), .B(n3257), .C(n65567), .Q(N2745) );
  OAI212 U6351 ( .A(n3253), .B(n3257), .C(n65568), .Q(N2744) );
  OAI212 U6353 ( .A(n3245), .B(n3258), .C(n65567), .Q(N2743) );
  OAI212 U6354 ( .A(n3247), .B(n3258), .C(n65568), .Q(N2742) );
  OAI212 U6355 ( .A(n3248), .B(n3258), .C(n65568), .Q(N2741) );
  OAI212 U6356 ( .A(n3249), .B(n3258), .C(n65567), .Q(N2740) );
  OAI212 U6357 ( .A(n3250), .B(n3258), .C(n65569), .Q(N2739) );
  OAI212 U6358 ( .A(n3251), .B(n3258), .C(n66568), .Q(N2738) );
  OAI212 U6359 ( .A(n3252), .B(n3258), .C(n65569), .Q(N2737) );
  OAI212 U6360 ( .A(n3253), .B(n3258), .C(n66568), .Q(N2736) );
  OAI212 U6362 ( .A(n3245), .B(n3259), .C(n65569), .Q(N2735) );
  OAI212 U6363 ( .A(n3247), .B(n3259), .C(n66568), .Q(N2734) );
  OAI212 U6364 ( .A(n3248), .B(n3259), .C(n65569), .Q(N2733) );
  OAI212 U6365 ( .A(n3249), .B(n3259), .C(n66568), .Q(N2732) );
  OAI212 U6366 ( .A(n3250), .B(n3259), .C(n65569), .Q(N2731) );
  OAI212 U6367 ( .A(n3251), .B(n3259), .C(n66568), .Q(N2730) );
  OAI212 U6368 ( .A(n3252), .B(n3259), .C(n65569), .Q(N2729) );
  OAI212 U6369 ( .A(n3253), .B(n3259), .C(n66568), .Q(N2728) );
  OAI212 U6371 ( .A(n3245), .B(n3260), .C(n65569), .Q(N2727) );
  OAI212 U6373 ( .A(n3247), .B(n3260), .C(n66568), .Q(N2726) );
  OAI212 U6375 ( .A(n3248), .B(n3260), .C(n65569), .Q(N2725) );
  OAI212 U6377 ( .A(n3249), .B(n3260), .C(n66568), .Q(N2724) );
  OAI212 U6379 ( .A(n3250), .B(n3260), .C(n65569), .Q(N2723) );
  OAI212 U6381 ( .A(n3251), .B(n3260), .C(n66568), .Q(N2722) );
  OAI212 U6383 ( .A(n3252), .B(n3260), .C(n65569), .Q(N2721) );
  OAI212 U6385 ( .A(n3253), .B(n3260), .C(n66568), .Q(N2720) );
  OAI222 U6458 ( .A(n65554), .B(n3331), .C(n3332), .D(n3333), .Q(n3329) );
  OAI212 U6459 ( .A(n3334), .B(n65592), .C(n65570), .Q(N2678) );
  OAI222 U6461 ( .A(n66528), .B(n3340), .C(n3330), .D(n3341), .Q(n3339) );
  OAI212 U6462 ( .A(n65553), .B(n3342), .C(n3343), .Q(n3338) );
  OAI222 U6464 ( .A(n3347), .B(n3348), .C(n3349), .D(n3350), .Q(n3346) );
  OAI222 U6465 ( .A(n3351), .B(n3352), .C(n3353), .D(n3354), .Q(n3345) );
  OAI222 U6468 ( .A(n66535), .B(n3360), .C(n66587), .D(n3361), .Q(n3359) );
  OAI212 U6469 ( .A(n3363), .B(n65591), .C(n65570), .Q(N2676) );
  OAI222 U6471 ( .A(n66471), .B(n66486), .C(n66535), .D(n3367), .Q(n3366) );
  OAI212 U6473 ( .A(n66587), .B(n3368), .C(n3369), .Q(n3365) );
  OAI222 U6475 ( .A(n3347), .B(n3372), .C(n3349), .D(n3373), .Q(n3371) );
  OAI222 U6476 ( .A(n3351), .B(n3374), .C(n3353), .D(n3375), .Q(n3370) );
  OAI212 U6481 ( .A(n3385), .B(n65590), .C(n65570), .Q(N2674) );
  OAI222 U6483 ( .A(n66535), .B(n3389), .C(n66590), .D(n3390), .Q(n3388) );
  OAI212 U6484 ( .A(n66587), .B(n3391), .C(n3392), .Q(n3387) );
  OAI222 U6486 ( .A(n3347), .B(n3395), .C(n3349), .D(n3396), .Q(n3394) );
  OAI222 U6487 ( .A(n3351), .B(n3397), .C(n3353), .D(n3398), .Q(n3393) );
  OAI222 U6490 ( .A(n65553), .B(n3331), .C(n3333), .D(n65554), .Q(n3400) );
  OAI212 U6491 ( .A(n3401), .B(n65592), .C(n65570), .Q(N2672) );
  OAI222 U6493 ( .A(n66529), .B(n3340), .C(n65553), .D(n3341), .Q(n3403) );
  OAI212 U6494 ( .A(n65554), .B(n3342), .C(n3404), .Q(n3402) );
  OAI222 U6496 ( .A(n3347), .B(n3407), .C(n3349), .D(n3408), .Q(n3406) );
  OAI222 U6499 ( .A(n3351), .B(n3411), .C(n3353), .D(n3412), .Q(n3405) );
  OAI222 U6504 ( .A(n66589), .B(n3419), .C(n3361), .D(n66592), .Q(n3418) );
  OAI212 U6505 ( .A(n3420), .B(n65591), .C(n65570), .Q(N2670) );
  OAI222 U6507 ( .A(n3367), .B(n66533), .C(n66589), .D(n3425), .Q(n3424) );
  OAI212 U6508 ( .A(n3368), .B(n66592), .C(n3426), .Q(n3423) );
  OAI222 U6510 ( .A(n3348), .B(n3429), .C(n3350), .D(n3430), .Q(n3428) );
  OAI222 U6511 ( .A(n3352), .B(n3431), .C(n3354), .D(n3432), .Q(n3427) );
  OAI212 U6515 ( .A(n3439), .B(n65590), .C(n65570), .Q(N2668) );
  OAI222 U6517 ( .A(n3389), .B(n66534), .C(n3390), .D(n66588), .Q(n3441) );
  OAI212 U6518 ( .A(n3391), .B(n66591), .C(n3442), .Q(n3440) );
  OAI222 U6520 ( .A(n3372), .B(n3429), .C(n3373), .D(n3430), .Q(n3444) );
  OAI222 U6521 ( .A(n3374), .B(n3431), .C(n3375), .D(n3432), .Q(n3443) );
  OAI222 U6524 ( .A(n3331), .B(n66591), .C(n3333), .D(n66588), .Q(n3446) );
  OAI212 U6525 ( .A(n3447), .B(n65592), .C(n65570), .Q(N2666) );
  OAI222 U6527 ( .A(n3340), .B(n66530), .C(n3341), .D(n66591), .Q(n3449) );
  OAI212 U6528 ( .A(n3342), .B(n66588), .C(n3450), .Q(n3448) );
  OAI222 U6530 ( .A(n3395), .B(n3429), .C(n3396), .D(n3430), .Q(n3452) );
  OAI222 U6531 ( .A(n3397), .B(n3431), .C(n3398), .D(n3432), .Q(n3451) );
  OAI222 U6534 ( .A(n66592), .B(n3419), .C(n66589), .D(n3361), .Q(n3454) );
  OAI212 U6537 ( .A(n3457), .B(n65591), .C(n65570), .Q(N2664) );
  OAI222 U6539 ( .A(n66532), .B(n3367), .C(n66592), .D(n3425), .Q(n3459) );
  OAI212 U6542 ( .A(n66589), .B(n3368), .C(n3462), .Q(n3458) );
  OAI222 U6544 ( .A(n3407), .B(n3429), .C(n3408), .D(n3430), .Q(n3464) );
  OAI222 U6549 ( .A(n3411), .B(n3431), .C(n3412), .D(n3432), .Q(n3463) );
  OAI212 U6558 ( .A(n3438), .B(n3332), .C(n3476), .Q(n3475) );
  OAI212 U6559 ( .A(n3477), .B(n65590), .C(n65570), .Q(N2662) );
  OAI222 U6561 ( .A(n66528), .B(n3389), .C(n3330), .D(n3390), .Q(n3479) );
  OAI212 U6562 ( .A(n3332), .B(n3391), .C(n3480), .Q(n3478) );
  OAI222 U6564 ( .A(n3348), .B(n3483), .C(n3350), .D(n3484), .Q(n3482) );
  OAI222 U6565 ( .A(n3352), .B(n3485), .C(n3354), .D(n3486), .Q(n3481) );
  OAI222 U6568 ( .A(n3331), .B(n66587), .C(n3333), .D(n66590), .Q(n3488) );
  OAI212 U6571 ( .A(n3491), .B(n65592), .C(n3335), .Q(N2660) );
  OAI222 U6573 ( .A(n3340), .B(n66527), .C(n3341), .D(n66587), .Q(n3493) );
  OAI212 U6576 ( .A(n3342), .B(n66590), .C(n3497), .Q(n3492) );
  OAI222 U6578 ( .A(n3372), .B(n3483), .C(n3373), .D(n3484), .Q(n3499) );
  OAI222 U6579 ( .A(n3374), .B(n3485), .C(n3375), .D(n3486), .Q(n3498) );
  OAI222 U6584 ( .A(n66587), .B(n3419), .C(n66590), .D(n3506), .Q(n3505) );
  OAI212 U6585 ( .A(n3507), .B(n65591), .C(n3335), .Q(N2658) );
  OAI222 U6587 ( .A(n66527), .B(n3510), .C(n66587), .D(n3425), .Q(n3509) );
  OAI212 U6588 ( .A(n66590), .B(n3511), .C(n3512), .Q(n3508) );
  OAI222 U6590 ( .A(n3395), .B(n3483), .C(n3396), .D(n3484), .Q(n3514) );
  OAI222 U6591 ( .A(n3397), .B(n3485), .C(n3398), .D(n3486), .Q(n3513) );
  OAI212 U6594 ( .A(n3438), .B(n65554), .C(n3476), .Q(n3516) );
  OAI212 U6595 ( .A(n3517), .B(n65590), .C(n3335), .Q(N2656) );
  OAI222 U6597 ( .A(n66529), .B(n3389), .C(n65553), .D(n3390), .Q(n3519) );
  OAI212 U6598 ( .A(n3330), .B(n3391), .C(n3520), .Q(n3518) );
  OAI222 U6600 ( .A(n3407), .B(n3483), .C(n3408), .D(n3484), .Q(n3522) );
  OAI222 U6603 ( .A(n3411), .B(n3485), .C(n3412), .D(n3486), .Q(n3521) );
  OAI212 U6609 ( .A(n3532), .B(n65592), .C(n3335), .Q(N2654) );
  OAI222 U6611 ( .A(n66532), .B(n66470), .C(n3341), .D(n66592), .Q(n3534) );
  OAI212 U6612 ( .A(n66589), .B(n3535), .C(n3536), .Q(n3533) );
  OAI222 U6614 ( .A(n3348), .B(n3539), .C(n3350), .D(n3540), .Q(n3538) );
  OAI222 U6615 ( .A(n3352), .B(n3541), .C(n3354), .D(n3542), .Q(n3537) );
  OAI222 U6618 ( .A(n3419), .B(n66591), .C(n66588), .D(n3506), .Q(n3544) );
  OAI212 U6619 ( .A(n3545), .B(n65591), .C(n3335), .Q(N2652) );
  OAI222 U6621 ( .A(n66530), .B(n3510), .C(n3425), .D(n66591), .Q(n3547) );
  OAI212 U6622 ( .A(n66588), .B(n3511), .C(n3548), .Q(n3546) );
  OAI222 U6624 ( .A(n3372), .B(n3539), .C(n3373), .D(n3540), .Q(n3550) );
  OAI222 U6625 ( .A(n3374), .B(n3541), .C(n3375), .D(n3542), .Q(n3549) );
  OAI222 U6628 ( .A(n3377), .B(n66591), .C(n3438), .D(n66588), .Q(n3552) );
  OAI212 U6629 ( .A(n3553), .B(n65592), .C(n3335), .Q(N2650) );
  OAI222 U6631 ( .A(n3389), .B(n66530), .C(n3390), .D(n66591), .Q(n3555) );
  OAI212 U6632 ( .A(n3391), .B(n66588), .C(n3556), .Q(n3554) );
  OAI222 U6634 ( .A(n3395), .B(n3539), .C(n3396), .D(n3540), .Q(n3558) );
  OAI222 U6635 ( .A(n3397), .B(n3541), .C(n3398), .D(n3542), .Q(n3557) );
  OAI212 U6641 ( .A(n3564), .B(n65591), .C(n3335), .Q(N2648) );
  OAI222 U6643 ( .A(n66533), .B(n66470), .C(n66589), .D(n3341), .Q(n3566) );
  OAI212 U6645 ( .A(n66592), .B(n3535), .C(n3568), .Q(n3565) );
  OAI222 U6647 ( .A(n3407), .B(n3539), .C(n3408), .D(n3540), .Q(n3570) );
  OAI222 U6652 ( .A(n3411), .B(n3541), .C(n3412), .D(n3542), .Q(n3569) );
  OAI222 U6660 ( .A(n65553), .B(n3419), .C(n3330), .D(n3506), .Q(n3573) );
  OAI212 U6661 ( .A(n3574), .B(n65592), .C(n65570), .Q(N2646) );
  OAI222 U6663 ( .A(n66529), .B(n3510), .C(n3332), .D(n3425), .Q(n3576) );
  OAI212 U6664 ( .A(n65554), .B(n3511), .C(n3577), .Q(n3575) );
  OAI222 U6666 ( .A(n3348), .B(n3580), .C(n3350), .D(n3581), .Q(n3579) );
  OAI222 U6667 ( .A(n3352), .B(n3582), .C(n3354), .D(n3583), .Q(n3578) );
  OAI222 U6670 ( .A(n66587), .B(n3377), .C(n66590), .D(n3438), .Q(n3585) );
  OAI212 U6673 ( .A(n3588), .B(n65590), .C(n65570), .Q(N2644) );
  OAI222 U6675 ( .A(n66527), .B(n3389), .C(n66587), .D(n3390), .Q(n3590) );
  OAI212 U6677 ( .A(n66590), .B(n3391), .C(n3591), .Q(n3589) );
  OAI222 U6679 ( .A(n3372), .B(n3580), .C(n3373), .D(n3581), .Q(n3593) );
  OAI222 U6680 ( .A(n3374), .B(n3582), .C(n3375), .D(n3583), .Q(n3592) );
  OAI212 U6686 ( .A(n3598), .B(n65591), .C(n65570), .Q(N2642) );
  OAI222 U6688 ( .A(n66587), .B(n3535), .C(n66351), .D(n3601), .Q(n3600) );
  OAI222 U6689 ( .A(n3581), .B(n3396), .C(n3580), .D(n3395), .Q(n3602) );
  OAI222 U6696 ( .A(n3583), .B(n3398), .C(n3582), .D(n3397), .Q(n3605) );
  OAI222 U6700 ( .A(n65554), .B(n3419), .C(n65553), .D(n3506), .Q(n3607) );
  OAI212 U6701 ( .A(n3608), .B(n65592), .C(n65570), .Q(N2640) );
  OAI222 U6703 ( .A(n66528), .B(n3510), .C(n65554), .D(n3425), .Q(n3610) );
  OAI212 U6706 ( .A(n65553), .B(n3511), .C(n3611), .Q(n3609) );
  OAI222 U6708 ( .A(n3407), .B(n3580), .C(n3408), .D(n3581), .Q(n3613) );
  OAI222 U6713 ( .A(n3411), .B(n3582), .C(n3412), .D(n3583), .Q(n3612) );
  OAI212 U6724 ( .A(n3625), .B(n65590), .C(n65570), .Q(N2638) );
  OAI222 U6726 ( .A(n3390), .B(n66592), .C(n66340), .D(n3601), .Q(n3627) );
  OAI222 U6727 ( .A(n3629), .B(n3350), .C(n3630), .D(n3348), .Q(n3628) );
  OAI222 U6733 ( .A(n3634), .B(n3354), .C(n3635), .D(n3352), .Q(n3633) );
  OAI212 U6742 ( .A(n3643), .B(n65590), .C(n65570), .Q(N2636) );
  OAI222 U6744 ( .A(n66591), .B(n3535), .C(n66338), .D(n3601), .Q(n3645) );
  OAI222 U6745 ( .A(n3629), .B(n3373), .C(n3630), .D(n3372), .Q(n3646) );
  OAI222 U6754 ( .A(n3634), .B(n3375), .C(n3635), .D(n3374), .Q(n3651) );
  OAI222 U6760 ( .A(n3419), .B(n66588), .C(n66591), .D(n3506), .Q(n3653) );
  OAI212 U6766 ( .A(n3657), .B(n65592), .C(n65570), .Q(N2634) );
  OAI222 U6768 ( .A(n66534), .B(n3510), .C(n3425), .D(n66588), .Q(n3659) );
  OAI212 U6773 ( .A(n66591), .B(n3511), .C(n3660), .Q(n3658) );
  OAI222 U6775 ( .A(n3395), .B(n3630), .C(n3396), .D(n3629), .Q(n3662) );
  OAI222 U6778 ( .A(n3397), .B(n3635), .C(n3398), .D(n3634), .Q(n3661) );
  OAI212 U6812 ( .A(n3678), .B(n65591), .C(n65570), .Q(N2632) );
  OAI212 U6814 ( .A(n3676), .B(n3655), .C(n66567), .Q(n3679) );
  OAI222 U6818 ( .A(n66589), .B(n3390), .C(n66335), .D(n3601), .Q(n3681) );
  OAI222 U6819 ( .A(n3629), .B(n3408), .C(n3630), .D(n3407), .Q(n3682) );
  OAI222 U6871 ( .A(n3634), .B(n3412), .C(n3635), .D(n3411), .Q(n3706) );
  IMUX23 U7368 ( .A(n3855), .B(n3856), .S(n65936), .Q(N1904) );
  ADD22 \add_168/U1_1_1  ( .A(N2012), .B(N2013), .CO(\add_168/carry [2]), .S(
        N2015) );
  ADD22 \add_168/U1_1_2  ( .A(N2011), .B(\add_168/carry [2]), .CO(
        \add_168/carry [3]), .S(N2016) );
  ADD22 \add_168/U1_1_3  ( .A(N2010), .B(\add_168/carry [3]), .CO(
        \add_168/carry [4]), .S(N2017) );
  ADD22 \add_168/U1_1_4  ( .A(N2009), .B(\add_168/carry [4]), .CO(
        \add_168/carry [5]), .S(N2018) );
  ADD22 \add_168/U1_1_5  ( .A(N2008), .B(\add_168/carry [5]), .CO(
        \add_168/carry [6]), .S(N2019) );
  ADD22 \add_168/U1_1_6  ( .A(N2007), .B(\add_168/carry [6]), .CO(
        \add_168/carry [7]), .S(N2020) );
  ADD22 \add_168/U1_1_7  ( .A(N2006), .B(\add_168/carry [7]), .CO(
        \add_168/carry [8]), .S(N2021) );
  ADD22 \add_168/U1_1_8  ( .A(N2005), .B(\add_168/carry [8]), .CO(
        \add_168/carry [9]), .S(N2022) );
  ADD22 \add_168/U1_1_9  ( .A(N2004), .B(\add_168/carry [9]), .CO(
        \add_168/carry [10]), .S(N2023) );
  ADD22 \add_168/U1_1_10  ( .A(N2003), .B(\add_168/carry [10]), .CO(
        \add_168/carry [11]), .S(N2024) );
  ADD22 \add_168/U1_1_11  ( .A(N2002), .B(\add_168/carry [11]), .CO(
        \add_168/carry [12]), .S(N2025) );
  ADD22 \add_168/U1_1_12  ( .A(N2001), .B(\add_168/carry [12]), .CO(
        \add_168/carry [13]), .S(N2026) );
  ADD22 \add_168/U1_1_13  ( .A(N2000), .B(\add_168/carry [13]), .CO(
        \add_168/carry [14]), .S(N2027) );
  ADD22 \add_168/U1_1_14  ( .A(N1999), .B(\add_168/carry [14]), .CO(
        \add_168/carry [15]), .S(N2028) );
  ADD22 \add_168/U1_1_15  ( .A(N1998), .B(\add_168/carry [15]), .CO(
        \add_168/carry [16]), .S(N2029) );
  ADD22 \add_168/U1_1_16  ( .A(N1997), .B(\add_168/carry [16]), .CO(
        \add_168/carry [17]), .S(N2030) );
  ADD22 \add_168/U1_1_17  ( .A(N1996), .B(\add_168/carry [17]), .CO(
        \add_168/carry [18]), .S(N2031) );
  ADD22 \add_168/U1_1_18  ( .A(N1995), .B(\add_168/carry [18]), .CO(
        \add_168/carry [19]), .S(N2032) );
  ADD22 \add_168/U1_1_19  ( .A(N1994), .B(\add_168/carry [19]), .CO(
        \add_168/carry [20]), .S(N2033) );
  ADD22 \add_168/U1_1_20  ( .A(N1993), .B(\add_168/carry [20]), .CO(
        \add_168/carry [21]), .S(N2034) );
  ADD22 \add_168/U1_1_21  ( .A(N1992), .B(\add_168/carry [21]), .CO(
        \add_168/carry [22]), .S(N2035) );
  ADD22 \add_168/U1_1_22  ( .A(N1991), .B(\add_168/carry [22]), .CO(
        \add_168/carry [23]), .S(N2036) );
  ADD22 \add_168/U1_1_23  ( .A(N1990), .B(\add_168/carry [23]), .CO(
        \add_168/carry [24]), .S(N2037) );
  ADD22 \add_168/U1_1_24  ( .A(N1989), .B(\add_168/carry [24]), .CO(
        \add_168/carry [25]), .S(N2038) );
  ADD22 \add_168/U1_1_25  ( .A(N1988), .B(\add_168/carry [25]), .CO(
        \add_168/carry [26]), .S(N2039) );
  ADD22 \add_168/U1_1_26  ( .A(N1987), .B(\add_168/carry [26]), .CO(
        \add_168/carry [27]), .S(N2040) );
  ADD22 \add_168/U1_1_27  ( .A(N1986), .B(\add_168/carry [27]), .CO(
        \add_168/carry [28]), .S(N2041) );
  ADD22 \add_168/U1_1_28  ( .A(N1985), .B(\add_168/carry [28]), .CO(
        \add_168/carry [29]), .S(N2042) );
  ADD22 \add_168/U1_1_29  ( .A(N1984), .B(\add_168/carry [29]), .CO(
        \add_168/carry [30]), .S(N2043) );
  ADD22 \add_168/U1_1_30  ( .A(N1983), .B(\add_168/carry [30]), .CO(
        \add_168/carry [31]), .S(N2044) );
  ADD22 \add_137/U1_1_1  ( .A(N1469), .B(N1470), .CO(\add_137/carry [2]), .S(
        N1472) );
  ADD22 \add_137/U1_1_2  ( .A(N1468), .B(\add_137/carry [2]), .CO(
        \add_137/carry [3]), .S(N1473) );
  ADD22 \add_137/U1_1_3  ( .A(N1467), .B(\add_137/carry [3]), .CO(
        \add_137/carry [4]), .S(N1474) );
  ADD22 \add_137/U1_1_4  ( .A(N1466), .B(\add_137/carry [4]), .CO(
        \add_137/carry [5]), .S(N1475) );
  ADD22 \add_137/U1_1_5  ( .A(N1465), .B(\add_137/carry [5]), .CO(
        \add_137/carry [6]), .S(N1476) );
  ADD22 \add_137/U1_1_6  ( .A(N1464), .B(\add_137/carry [6]), .CO(
        \add_137/carry [7]), .S(N1477) );
  ADD22 \add_137/U1_1_7  ( .A(N1463), .B(\add_137/carry [7]), .CO(
        \add_137/carry [8]), .S(N1478) );
  ADD22 \add_137/U1_1_8  ( .A(N1462), .B(\add_137/carry [8]), .CO(
        \add_137/carry [9]), .S(N1479) );
  ADD22 \add_137/U1_1_9  ( .A(N1461), .B(\add_137/carry [9]), .CO(
        \add_137/carry [10]), .S(N1480) );
  ADD22 \add_137/U1_1_10  ( .A(N1460), .B(\add_137/carry [10]), .CO(
        \add_137/carry [11]), .S(N1481) );
  ADD22 \add_137/U1_1_11  ( .A(N1459), .B(\add_137/carry [11]), .CO(
        \add_137/carry [12]), .S(N1482) );
  ADD22 \add_137/U1_1_12  ( .A(N1458), .B(\add_137/carry [12]), .CO(
        \add_137/carry [13]), .S(N1483) );
  ADD22 \add_137/U1_1_13  ( .A(N1457), .B(\add_137/carry [13]), .CO(
        \add_137/carry [14]), .S(N1484) );
  ADD22 \add_137/U1_1_14  ( .A(N1456), .B(\add_137/carry [14]), .CO(
        \add_137/carry [15]), .S(N1485) );
  ADD22 \add_137/U1_1_15  ( .A(N1455), .B(\add_137/carry [15]), .CO(
        \add_137/carry [16]), .S(N1486) );
  ADD22 \add_137/U1_1_16  ( .A(N1454), .B(\add_137/carry [16]), .CO(
        \add_137/carry [17]), .S(N1487) );
  ADD22 \add_137/U1_1_17  ( .A(N1453), .B(\add_137/carry [17]), .CO(
        \add_137/carry [18]), .S(N1488) );
  ADD22 \add_137/U1_1_18  ( .A(N1452), .B(\add_137/carry [18]), .CO(
        \add_137/carry [19]), .S(N1489) );
  ADD22 \add_137/U1_1_19  ( .A(N1451), .B(\add_137/carry [19]), .CO(
        \add_137/carry [20]), .S(N1490) );
  ADD22 \add_137/U1_1_20  ( .A(N1450), .B(\add_137/carry [20]), .CO(
        \add_137/carry [21]), .S(N1491) );
  ADD22 \add_137/U1_1_21  ( .A(N1449), .B(\add_137/carry [21]), .CO(
        \add_137/carry [22]), .S(N1492) );
  ADD22 \add_137/U1_1_22  ( .A(N1448), .B(\add_137/carry [22]), .CO(
        \add_137/carry [23]), .S(N1493) );
  ADD22 \add_137/U1_1_23  ( .A(N1447), .B(\add_137/carry [23]), .CO(
        \add_137/carry [24]), .S(N1494) );
  ADD22 \add_137/U1_1_24  ( .A(N1446), .B(\add_137/carry [24]), .CO(
        \add_137/carry [25]), .S(N1495) );
  ADD22 \add_137/U1_1_25  ( .A(N1445), .B(\add_137/carry [25]), .CO(
        \add_137/carry [26]), .S(N1496) );
  ADD22 \add_137/U1_1_26  ( .A(N1444), .B(\add_137/carry [26]), .CO(
        \add_137/carry [27]), .S(N1497) );
  ADD22 \add_137/U1_1_27  ( .A(N1443), .B(\add_137/carry [27]), .CO(
        \add_137/carry [28]), .S(N1498) );
  ADD22 \add_137/U1_1_28  ( .A(N1442), .B(\add_137/carry [28]), .CO(
        \add_137/carry [29]), .S(N1499) );
  ADD22 \add_137/U1_1_29  ( .A(N1441), .B(\add_137/carry [29]), .CO(
        \add_137/carry [30]), .S(N1500) );
  ADD22 \add_137/U1_1_30  ( .A(N1440), .B(\add_137/carry [30]), .CO(
        \add_137/carry [31]), .S(N1501) );
  DF3 \G_play_reg[3]  ( .D(G[3]), .C(CLK), .QN(n1680) );
  DLPQ3 \m_reg[0]  ( .SN(n807), .D(N2849), .GN(n66393), .Q(N3200) );
  DF3 \C4_OUT_reg[0]  ( .D(n65436), .C(CLK), .Q(C4_OUT[0]), .QN(n1682) );
  DLPQ3 \next_state_reg[0]  ( .SN(n807), .D(N2630), .GN(n66566), .Q(
        next_state[0]) );
  DFC3 \state_reg[0]  ( .D(next_state[0]), .C(CLK), .RN(NRST), .Q(state[0]), 
        .QN(n1654) );
  DLPQ3 \next_state_reg[1]  ( .SN(n807), .D(n65587), .GN(n66566), .Q(
        next_state[1]) );
  DFC3 \state_reg[1]  ( .D(next_state[1]), .C(CLK), .RN(NRST), .Q(state[1]) );
  DLPQ3 \GFill_reg[0][0]  ( .SN(n807), .D(n65588), .GN(n66227), .Q(
        \GFill[0][0] ) );
  DLPQ3 \GFill_reg[1][0]  ( .SN(n807), .D(n65588), .GN(n66228), .Q(
        \GFill[1][0] ) );
  DLPQ3 \GFill_reg[2][0]  ( .SN(n807), .D(n65589), .GN(n66229), .Q(
        \GFill[2][0] ) );
  DLPQ3 \GFill_reg[3][0]  ( .SN(n807), .D(n65588), .GN(n66230), .Q(
        \GFill[3][0] ) );
  DLPQ3 \GFill_reg[4][0]  ( .SN(n807), .D(n65588), .GN(n66231), .Q(
        \GFill[4][0] ) );
  DLPQ3 \GFill_reg[5][0]  ( .SN(n807), .D(n65587), .GN(n66232), .Q(
        \GFill[5][0] ) );
  DLPQ3 \GFill_reg[6][0]  ( .SN(n807), .D(n65586), .GN(n66233), .Q(
        \GFill[6][0] ) );
  DLPQ3 \GFill_reg[7][0]  ( .SN(n807), .D(n65587), .GN(n66234), .Q(
        \GFill[7][0] ) );
  DLPQ3 \GFill_reg[8][0]  ( .SN(n807), .D(n65586), .GN(n66219), .Q(
        \GFill[8][0] ) );
  DLPQ3 \GFill_reg[9][0]  ( .SN(n807), .D(n65587), .GN(n66220), .Q(
        \GFill[9][0] ) );
  DLPQ3 \GFill_reg[10][0]  ( .SN(n807), .D(n65586), .GN(n66221), .Q(
        \GFill[10][0] ) );
  DLPQ3 \GFill_reg[11][0]  ( .SN(n807), .D(n65586), .GN(n66222), .Q(
        \GFill[11][0] ) );
  DLPQ3 \GFill_reg[12][0]  ( .SN(n807), .D(n65589), .GN(n66223), .Q(
        \GFill[12][0] ) );
  DLPQ3 \GFill_reg[13][0]  ( .SN(n807), .D(n65588), .GN(n66224), .Q(
        \GFill[13][0] ) );
  DLPQ3 \GFill_reg[14][0]  ( .SN(n807), .D(n65589), .GN(n66225), .Q(
        \GFill[14][0] ) );
  DLPQ3 \GFill_reg[15][0]  ( .SN(n807), .D(n65588), .GN(n66226), .Q(
        \GFill[15][0] ) );
  DLPQ3 \GFill_reg[16][0]  ( .SN(n807), .D(n65587), .GN(n66211), .Q(
        \GFill[16][0] ) );
  DLPQ3 \GFill_reg[17][0]  ( .SN(n807), .D(n65587), .GN(n66212), .Q(
        \GFill[17][0] ) );
  DLPQ3 \GFill_reg[18][0]  ( .SN(n807), .D(n65586), .GN(n66213), .Q(
        \GFill[18][0] ) );
  DLPQ3 \GFill_reg[19][0]  ( .SN(n807), .D(n65586), .GN(n66214), .Q(
        \GFill[19][0] ) );
  DLPQ3 \GFill_reg[20][0]  ( .SN(n807), .D(n65586), .GN(n66215), .Q(
        \GFill[20][0] ) );
  DLPQ3 \GFill_reg[21][0]  ( .SN(n807), .D(n65587), .GN(n66216), .Q(
        \GFill[21][0] ) );
  DLPQ3 \GFill_reg[22][0]  ( .SN(n807), .D(n65589), .GN(n66217), .Q(
        \GFill[22][0] ) );
  DLPQ3 \GFill_reg[23][0]  ( .SN(n807), .D(n65586), .GN(n66218), .Q(
        \GFill[23][0] ) );
  DLPQ3 \GFill_reg[24][0]  ( .SN(n807), .D(n65588), .GN(n66203), .Q(
        \GFill[24][0] ) );
  DLPQ3 \GFill_reg[25][0]  ( .SN(n807), .D(n65587), .GN(n66204), .Q(
        \GFill[25][0] ) );
  DLPQ3 \GFill_reg[26][0]  ( .SN(n807), .D(n65588), .GN(n66205), .Q(
        \GFill[26][0] ) );
  DLPQ3 \GFill_reg[27][0]  ( .SN(n807), .D(n65586), .GN(n66206), .Q(
        \GFill[27][0] ) );
  DLPQ3 \GFill_reg[28][0]  ( .SN(n807), .D(n65588), .GN(n66207), .Q(
        \GFill[28][0] ) );
  DLPQ3 \GFill_reg[29][0]  ( .SN(n807), .D(N2631), .GN(n66208), .Q(
        \GFill[29][0] ) );
  DLPQ3 \GFill_reg[30][0]  ( .SN(n807), .D(n65586), .GN(n66209), .Q(
        \GFill[30][0] ) );
  DLPQ3 \GFill_reg[31][0]  ( .SN(n807), .D(n65586), .GN(n66210), .Q(
        \GFill[31][0] ) );
  DLPQ3 \GFill_reg[32][0]  ( .SN(n807), .D(n65589), .GN(n66195), .Q(
        \GFill[32][0] ) );
  DLPQ3 \GFill_reg[33][0]  ( .SN(n807), .D(n65588), .GN(n66196), .Q(
        \GFill[33][0] ) );
  DLPQ3 \GFill_reg[34][0]  ( .SN(n807), .D(n65588), .GN(n66197), .Q(
        \GFill[34][0] ) );
  DLPQ3 \GFill_reg[35][0]  ( .SN(n807), .D(n65587), .GN(n66198), .Q(
        \GFill[35][0] ) );
  DLPQ3 \GFill_reg[36][0]  ( .SN(n807), .D(n65588), .GN(n66199), .Q(
        \GFill[36][0] ) );
  DLPQ3 \GFill_reg[37][0]  ( .SN(n807), .D(n65587), .GN(n66200), .Q(
        \GFill[37][0] ) );
  DLPQ3 \GFill_reg[38][0]  ( .SN(n807), .D(n65589), .GN(n66201), .Q(
        \GFill[38][0] ) );
  DLPQ3 \GFill_reg[39][0]  ( .SN(n807), .D(n65586), .GN(n66202), .Q(
        \GFill[39][0] ) );
  DLPQ3 \GFill_reg[40][0]  ( .SN(n807), .D(n65589), .GN(n66187), .Q(
        \GFill[40][0] ) );
  DLPQ3 \GFill_reg[41][0]  ( .SN(n807), .D(n65589), .GN(n66188), .Q(
        \GFill[41][0] ) );
  DLPQ3 \GFill_reg[42][0]  ( .SN(n807), .D(N2631), .GN(n66189), .Q(
        \GFill[42][0] ) );
  DLPQ3 \GFill_reg[43][0]  ( .SN(n807), .D(N2631), .GN(n66190), .Q(
        \GFill[43][0] ) );
  DLPQ3 \GFill_reg[44][0]  ( .SN(n807), .D(n65586), .GN(n66191), .Q(
        \GFill[44][0] ) );
  DLPQ3 \GFill_reg[45][0]  ( .SN(n807), .D(n65586), .GN(n66192), .Q(
        \GFill[45][0] ) );
  DLPQ3 \GFill_reg[46][0]  ( .SN(n807), .D(n65586), .GN(n66193), .Q(
        \GFill[46][0] ) );
  DLPQ3 \GFill_reg[47][0]  ( .SN(n807), .D(n65586), .GN(n66194), .Q(
        \GFill[47][0] ) );
  DLPQ3 \GFill_reg[48][0]  ( .SN(n807), .D(n65586), .GN(n66179), .Q(
        \GFill[48][0] ) );
  DLPQ3 \GFill_reg[49][0]  ( .SN(n807), .D(n65589), .GN(n66180), .Q(
        \GFill[49][0] ) );
  DLPQ3 \GFill_reg[50][0]  ( .SN(n807), .D(n65588), .GN(n66181), .Q(
        \GFill[50][0] ) );
  DLPQ3 \GFill_reg[51][0]  ( .SN(n807), .D(n65587), .GN(n66182), .Q(
        \GFill[51][0] ) );
  DLPQ3 \GFill_reg[52][0]  ( .SN(n807), .D(n65586), .GN(n66183), .Q(
        \GFill[52][0] ) );
  DLPQ3 \GFill_reg[53][0]  ( .SN(n807), .D(n65589), .GN(n66184), .Q(
        \GFill[53][0] ) );
  DLPQ3 \GFill_reg[54][0]  ( .SN(n807), .D(n65589), .GN(n66185), .Q(
        \GFill[54][0] ) );
  DLPQ3 \GFill_reg[55][0]  ( .SN(n807), .D(n65589), .GN(n66186), .Q(
        \GFill[55][0] ) );
  DLPQ3 \GFill_reg[56][0]  ( .SN(n807), .D(n65588), .GN(n66171), .Q(
        \GFill[56][0] ) );
  DLPQ3 \GFill_reg[57][0]  ( .SN(n807), .D(n65587), .GN(n66172), .Q(
        \GFill[57][0] ) );
  DLPQ3 \GFill_reg[58][0]  ( .SN(n807), .D(N2631), .GN(n66173), .Q(
        \GFill[58][0] ) );
  DLPQ3 \GFill_reg[59][0]  ( .SN(n807), .D(n65589), .GN(n66174), .Q(
        \GFill[59][0] ) );
  DLPQ3 \GFill_reg[60][0]  ( .SN(n807), .D(n65589), .GN(n66175), .Q(
        \GFill[60][0] ) );
  DLPQ3 \GFill_reg[61][0]  ( .SN(n807), .D(n65588), .GN(n66176), .Q(
        \GFill[61][0] ) );
  DLPQ3 \GFill_reg[62][0]  ( .SN(n807), .D(n65588), .GN(n66177), .Q(
        \GFill[62][0] ) );
  DLPQ3 \GFill_reg[63][0]  ( .SN(n807), .D(n65588), .GN(n66178), .Q(
        \GFill[63][0] ) );
  DLPQ3 \Col_Fill_reg[0][31]  ( .SN(n807), .D(n66466), .GN(n66375), .Q(
        \Col_Fill[0][31] ) );
  DLPQ3 \Col_Fill_reg[1][31]  ( .SN(n807), .D(n66466), .GN(n66376), .Q(
        \Col_Fill[1][31] ) );
  DLPQ3 \m_reg[3]  ( .SN(n807), .D(n66384), .GN(n66393), .Q(m[3]) );
  DLPQ3 \m_reg[2]  ( .SN(n807), .D(n66432), .GN(n66393), .Q(m[2]) );
  DLPQ3 \m_reg[1]  ( .SN(n807), .D(n66433), .GN(n66393), .Q(m[1]) );
  DLPQ3 \OFill_reg[63][0]  ( .SN(n807), .D(n65589), .GN(n66251), .Q(
        \OFill[63][0] ) );
  DLPQ3 \OFill_reg[62][0]  ( .SN(n807), .D(n65589), .GN(n66250), .Q(
        \OFill[62][0] ) );
  DLPQ3 \OFill_reg[61][0]  ( .SN(n807), .D(n65588), .GN(n66249), .Q(
        \OFill[61][0] ) );
  DLPQ3 \OFill_reg[60][0]  ( .SN(n807), .D(n65589), .GN(n66248), .Q(
        \OFill[60][0] ) );
  DLPQ3 \OFill_reg[59][0]  ( .SN(n807), .D(n65589), .GN(n66247), .Q(
        \OFill[59][0] ) );
  DLPQ3 \OFill_reg[58][0]  ( .SN(n807), .D(n65587), .GN(n66246), .Q(
        \OFill[58][0] ) );
  DLPQ3 \OFill_reg[57][0]  ( .SN(n807), .D(n65588), .GN(n66245), .Q(
        \OFill[57][0] ) );
  DLPQ3 \OFill_reg[56][0]  ( .SN(n807), .D(n65589), .GN(n66244), .Q(
        \OFill[56][0] ) );
  DLPQ3 \OFill_reg[55][0]  ( .SN(n807), .D(n65586), .GN(n66259), .Q(
        \OFill[55][0] ) );
  DLPQ3 \OFill_reg[54][0]  ( .SN(n807), .D(n65587), .GN(n66258), .Q(
        \OFill[54][0] ) );
  DLPQ3 \OFill_reg[53][0]  ( .SN(n807), .D(n65586), .GN(n66257), .Q(
        \OFill[53][0] ) );
  DLPQ3 \OFill_reg[52][0]  ( .SN(n807), .D(n65589), .GN(n66256), .Q(
        \OFill[52][0] ) );
  DLPQ3 \OFill_reg[51][0]  ( .SN(n807), .D(n65589), .GN(n66255), .Q(
        \OFill[51][0] ) );
  DLPQ3 \OFill_reg[50][0]  ( .SN(n807), .D(n65587), .GN(n66254), .Q(
        \OFill[50][0] ) );
  DLPQ3 \OFill_reg[49][0]  ( .SN(n807), .D(N2631), .GN(n66253), .Q(
        \OFill[49][0] ) );
  DLPQ3 \OFill_reg[48][0]  ( .SN(n807), .D(n65588), .GN(n66252), .Q(
        \OFill[48][0] ) );
  DLPQ3 \OFill_reg[47][0]  ( .SN(n807), .D(n65586), .GN(n66267), .Q(
        \OFill[47][0] ) );
  DLPQ3 \OFill_reg[46][0]  ( .SN(n807), .D(n65586), .GN(n66266), .Q(
        \OFill[46][0] ) );
  DLPQ3 \OFill_reg[45][0]  ( .SN(n807), .D(n65589), .GN(n66265), .Q(
        \OFill[45][0] ) );
  DLPQ3 \OFill_reg[44][0]  ( .SN(n807), .D(n65586), .GN(n66264), .Q(
        \OFill[44][0] ) );
  DLPQ3 \OFill_reg[43][0]  ( .SN(n807), .D(n65587), .GN(n66263), .Q(
        \OFill[43][0] ) );
  DLPQ3 \OFill_reg[42][0]  ( .SN(n807), .D(n65587), .GN(n66262), .Q(
        \OFill[42][0] ) );
  DLPQ3 \OFill_reg[41][0]  ( .SN(n807), .D(n65586), .GN(n66261), .Q(
        \OFill[41][0] ) );
  DLPQ3 \OFill_reg[40][0]  ( .SN(n807), .D(N2631), .GN(n66260), .Q(
        \OFill[40][0] ) );
  DLPQ3 \OFill_reg[39][0]  ( .SN(n807), .D(n65588), .GN(n66275), .Q(
        \OFill[39][0] ) );
  DLPQ3 \OFill_reg[38][0]  ( .SN(n807), .D(n65587), .GN(n66274), .Q(
        \OFill[38][0] ) );
  DLPQ3 \OFill_reg[37][0]  ( .SN(n807), .D(n65587), .GN(n66273), .Q(
        \OFill[37][0] ) );
  DLPQ3 \OFill_reg[36][0]  ( .SN(n807), .D(n65587), .GN(n66272), .Q(
        \OFill[36][0] ) );
  DLPQ3 \OFill_reg[35][0]  ( .SN(n807), .D(n65587), .GN(n66271), .Q(
        \OFill[35][0] ) );
  DLPQ3 \OFill_reg[34][0]  ( .SN(n807), .D(n65587), .GN(n66270), .Q(
        \OFill[34][0] ) );
  DLPQ3 \OFill_reg[33][0]  ( .SN(n807), .D(n65588), .GN(n66269), .Q(
        \OFill[33][0] ) );
  DLPQ3 \OFill_reg[32][0]  ( .SN(n807), .D(n65588), .GN(n66268), .Q(
        \OFill[32][0] ) );
  DLPQ3 \OFill_reg[31][0]  ( .SN(n807), .D(n65588), .GN(n66283), .Q(
        \OFill[31][0] ) );
  DLPQ3 \OFill_reg[30][0]  ( .SN(n807), .D(n65588), .GN(n66282), .Q(
        \OFill[30][0] ) );
  DLPQ3 \OFill_reg[29][0]  ( .SN(n807), .D(n65588), .GN(n66281), .Q(
        \OFill[29][0] ) );
  DLPQ3 \OFill_reg[28][0]  ( .SN(n807), .D(n65589), .GN(n66280), .Q(
        \OFill[28][0] ) );
  DLPQ3 \OFill_reg[27][0]  ( .SN(n807), .D(n65589), .GN(n66279), .Q(
        \OFill[27][0] ) );
  DLPQ3 \OFill_reg[26][0]  ( .SN(n807), .D(n65589), .GN(n66278), .Q(
        \OFill[26][0] ) );
  DLPQ3 \OFill_reg[25][0]  ( .SN(n807), .D(n65589), .GN(n66277), .Q(
        \OFill[25][0] ) );
  DLPQ3 \OFill_reg[24][0]  ( .SN(n807), .D(n65589), .GN(n66276), .Q(
        \OFill[24][0] ) );
  DLPQ3 \OFill_reg[23][0]  ( .SN(n807), .D(n65587), .GN(n66291), .Q(
        \OFill[23][0] ) );
  DLPQ3 \OFill_reg[22][0]  ( .SN(n807), .D(n65587), .GN(n66290), .Q(
        \OFill[22][0] ) );
  DLPQ3 \OFill_reg[21][0]  ( .SN(n807), .D(n65586), .GN(n66289), .Q(
        \OFill[21][0] ) );
  DLPQ3 \OFill_reg[20][0]  ( .SN(n807), .D(n65588), .GN(n66288), .Q(
        \OFill[20][0] ) );
  DLPQ3 \OFill_reg[19][0]  ( .SN(n807), .D(n65589), .GN(n66287), .Q(
        \OFill[19][0] ) );
  DLPQ3 \OFill_reg[18][0]  ( .SN(n807), .D(n65587), .GN(n66286), .Q(
        \OFill[18][0] ) );
  DLPQ3 \OFill_reg[17][0]  ( .SN(n807), .D(n65587), .GN(n66285), .Q(
        \OFill[17][0] ) );
  DLPQ3 \OFill_reg[16][0]  ( .SN(n807), .D(n65586), .GN(n66284), .Q(
        \OFill[16][0] ) );
  DLPQ3 \OFill_reg[15][0]  ( .SN(n807), .D(n65587), .GN(n66299), .Q(
        \OFill[15][0] ) );
  DLPQ3 \OFill_reg[14][0]  ( .SN(n807), .D(n65588), .GN(n66298), .Q(
        \OFill[14][0] ) );
  DLPQ3 \OFill_reg[13][0]  ( .SN(n807), .D(n65588), .GN(n66297), .Q(
        \OFill[13][0] ) );
  DLPQ3 \OFill_reg[12][0]  ( .SN(n807), .D(n65589), .GN(n66296), .Q(
        \OFill[12][0] ) );
  DLPQ3 \OFill_reg[11][0]  ( .SN(n807), .D(n65588), .GN(n66295), .Q(
        \OFill[11][0] ) );
  DLPQ3 \OFill_reg[10][0]  ( .SN(n807), .D(n65586), .GN(n66294), .Q(
        \OFill[10][0] ) );
  DLPQ3 \OFill_reg[9][0]  ( .SN(n807), .D(n65586), .GN(n66293), .Q(
        \OFill[9][0] ) );
  DLPQ3 \OFill_reg[8][0]  ( .SN(n807), .D(n65587), .GN(n66292), .Q(
        \OFill[8][0] ) );
  DLPQ3 \OFill_reg[7][0]  ( .SN(n807), .D(n65589), .GN(n66307), .Q(
        \OFill[7][0] ) );
  DLPQ3 \OFill_reg[6][0]  ( .SN(n807), .D(n65586), .GN(n66306), .Q(
        \OFill[6][0] ) );
  DLPQ3 \OFill_reg[5][0]  ( .SN(n807), .D(n65586), .GN(n66305), .Q(
        \OFill[5][0] ) );
  DLPQ3 \OFill_reg[4][0]  ( .SN(n807), .D(n65587), .GN(n66304), .Q(
        \OFill[4][0] ) );
  DLPQ3 \OFill_reg[3][0]  ( .SN(n807), .D(N2631), .GN(n66303), .Q(
        \OFill[3][0] ) );
  DLPQ3 \OFill_reg[2][0]  ( .SN(n807), .D(N2631), .GN(n66302), .Q(
        \OFill[2][0] ) );
  DLPQ3 \OFill_reg[1][0]  ( .SN(n807), .D(N2631), .GN(n66301), .Q(
        \OFill[1][0] ) );
  DLPQ3 \OFill_reg[0][0]  ( .SN(n807), .D(N2631), .GN(n66300), .Q(
        \OFill[0][0] ) );
  DLPQ3 \Col_Fill_reg[7][31]  ( .SN(n807), .D(n66466), .GN(n66382), .Q(
        \Col_Fill[7][31] ) );
  DLPQ3 \Col_Fill_reg[6][31]  ( .SN(n807), .D(n66466), .GN(n66381), .Q(
        \Col_Fill[6][31] ) );
  DLPQ3 \Col_Fill_reg[5][31]  ( .SN(n807), .D(n66466), .GN(n65561), .Q(
        \Col_Fill[5][31] ) );
  DLPQ3 \Col_Fill_reg[4][31]  ( .SN(n807), .D(n66466), .GN(n66379), .Q(
        \Col_Fill[4][31] ) );
  DLPQ3 \Col_Fill_reg[3][31]  ( .SN(n807), .D(n66466), .GN(n66378), .Q(
        \Col_Fill[3][31] ) );
  DLPQ3 \Col_Fill_reg[2][31]  ( .SN(n807), .D(n66466), .GN(n66377), .Q(
        \Col_Fill[2][31] ) );
  DLPQ3 \Col_Fill_reg[1][30]  ( .SN(n807), .D(n66465), .GN(n66376), .Q(
        \Col_Fill[1][30] ) );
  DLPQ3 \Col_Fill_reg[7][0]  ( .SN(n807), .D(n66435), .GN(n66382), .Q(
        \Col_Fill[7][0] ) );
  DLPQ3 \Col_Fill_reg[6][0]  ( .SN(n807), .D(n66435), .GN(n65562), .Q(
        \Col_Fill[6][0] ) );
  DLPQ3 \Col_Fill_reg[5][0]  ( .SN(n807), .D(n66435), .GN(n65561), .Q(
        \Col_Fill[5][0] ) );
  DLPQ3 \Col_Fill_reg[4][0]  ( .SN(n807), .D(n66435), .GN(n66379), .Q(
        \Col_Fill[4][0] ) );
  DLPQ3 \Col_Fill_reg[3][0]  ( .SN(n807), .D(n66435), .GN(n65559), .Q(
        \Col_Fill[3][0] ) );
  DLPQ3 \Col_Fill_reg[2][0]  ( .SN(n807), .D(n66435), .GN(n66377), .Q(
        \Col_Fill[2][0] ) );
  DLPQ3 \Col_Fill_reg[1][0]  ( .SN(n807), .D(n66435), .GN(n66376), .Q(
        \Col_Fill[1][0] ) );
  DLPQ3 \Col_Fill_reg[0][0]  ( .SN(n807), .D(n66435), .GN(n66375), .Q(
        \Col_Fill[0][0] ) );
  DLPQ3 \Col_Fill_reg[7][1]  ( .SN(n807), .D(n66436), .GN(n66382), .Q(
        \Col_Fill[7][1] ) );
  DLPQ3 \Col_Fill_reg[6][1]  ( .SN(n807), .D(n66436), .GN(n66381), .Q(
        \Col_Fill[6][1] ) );
  DLPQ3 \Col_Fill_reg[5][1]  ( .SN(n807), .D(n66436), .GN(n65561), .Q(
        \Col_Fill[5][1] ) );
  DLPQ3 \Col_Fill_reg[4][1]  ( .SN(n807), .D(n66436), .GN(n66379), .Q(
        \Col_Fill[4][1] ) );
  DLPQ3 \Col_Fill_reg[3][1]  ( .SN(n807), .D(n66436), .GN(n66378), .Q(
        \Col_Fill[3][1] ) );
  DLPQ3 \Col_Fill_reg[2][1]  ( .SN(n807), .D(n66436), .GN(n66377), .Q(
        \Col_Fill[2][1] ) );
  DLPQ3 \Col_Fill_reg[1][1]  ( .SN(n807), .D(n66436), .GN(n66376), .Q(
        \Col_Fill[1][1] ) );
  DLPQ3 \Col_Fill_reg[0][1]  ( .SN(n807), .D(n66436), .GN(n66375), .Q(
        \Col_Fill[0][1] ) );
  DLPQ3 \Col_Fill_reg[7][2]  ( .SN(n807), .D(n66437), .GN(n66382), .Q(
        \Col_Fill[7][2] ) );
  DLPQ3 \Col_Fill_reg[6][2]  ( .SN(n807), .D(n66437), .GN(n66381), .Q(
        \Col_Fill[6][2] ) );
  DLPQ3 \Col_Fill_reg[5][2]  ( .SN(n807), .D(n66437), .GN(n65561), .Q(
        \Col_Fill[5][2] ) );
  DLPQ3 \Col_Fill_reg[4][2]  ( .SN(n807), .D(n66437), .GN(n66379), .Q(
        \Col_Fill[4][2] ) );
  DLPQ3 \Col_Fill_reg[3][2]  ( .SN(n807), .D(n66437), .GN(n66378), .Q(
        \Col_Fill[3][2] ) );
  DLPQ3 \Col_Fill_reg[2][2]  ( .SN(n807), .D(n66437), .GN(n66377), .Q(
        \Col_Fill[2][2] ) );
  DLPQ3 \Col_Fill_reg[1][2]  ( .SN(n807), .D(n66437), .GN(n66376), .Q(
        \Col_Fill[1][2] ) );
  DLPQ3 \Col_Fill_reg[0][2]  ( .SN(n807), .D(n66437), .GN(n66375), .Q(
        \Col_Fill[0][2] ) );
  DLPQ3 \Col_Fill_reg[7][3]  ( .SN(n807), .D(n66438), .GN(n66382), .Q(
        \Col_Fill[7][3] ) );
  DLPQ3 \Col_Fill_reg[6][3]  ( .SN(n807), .D(n66438), .GN(n66381), .Q(
        \Col_Fill[6][3] ) );
  DLPQ3 \Col_Fill_reg[5][3]  ( .SN(n807), .D(n66438), .GN(n66380), .Q(
        \Col_Fill[5][3] ) );
  DLPQ3 \Col_Fill_reg[4][3]  ( .SN(n807), .D(n66438), .GN(n66379), .Q(
        \Col_Fill[4][3] ) );
  DLPQ3 \Col_Fill_reg[3][3]  ( .SN(n807), .D(n66438), .GN(n66378), .Q(
        \Col_Fill[3][3] ) );
  DLPQ3 \Col_Fill_reg[2][3]  ( .SN(n807), .D(n66438), .GN(n66377), .Q(
        \Col_Fill[2][3] ) );
  DLPQ3 \Col_Fill_reg[1][3]  ( .SN(n807), .D(n66438), .GN(n65557), .Q(
        \Col_Fill[1][3] ) );
  DLPQ3 \Col_Fill_reg[0][3]  ( .SN(n807), .D(n66438), .GN(n66375), .Q(
        \Col_Fill[0][3] ) );
  DLPQ3 \Col_Fill_reg[7][4]  ( .SN(n807), .D(n66439), .GN(n65563), .Q(
        \Col_Fill[7][4] ) );
  DLPQ3 \Col_Fill_reg[6][4]  ( .SN(n807), .D(n66439), .GN(n65562), .Q(
        \Col_Fill[6][4] ) );
  DLPQ3 \Col_Fill_reg[5][4]  ( .SN(n807), .D(n66439), .GN(n65561), .Q(
        \Col_Fill[5][4] ) );
  DLPQ3 \Col_Fill_reg[4][4]  ( .SN(n807), .D(n66439), .GN(n65560), .Q(
        \Col_Fill[4][4] ) );
  DLPQ3 \Col_Fill_reg[3][4]  ( .SN(n807), .D(n66439), .GN(n65559), .Q(
        \Col_Fill[3][4] ) );
  DLPQ3 \Col_Fill_reg[2][4]  ( .SN(n807), .D(n66439), .GN(n65558), .Q(
        \Col_Fill[2][4] ) );
  DLPQ3 \Col_Fill_reg[1][4]  ( .SN(n807), .D(n66439), .GN(n65557), .Q(
        \Col_Fill[1][4] ) );
  DLPQ3 \Col_Fill_reg[0][4]  ( .SN(n807), .D(n66439), .GN(n65556), .Q(
        \Col_Fill[0][4] ) );
  DLPQ3 \Col_Fill_reg[7][5]  ( .SN(n807), .D(n66440), .GN(n65563), .Q(
        \Col_Fill[7][5] ) );
  DLPQ3 \Col_Fill_reg[6][5]  ( .SN(n807), .D(n66440), .GN(n66381), .Q(
        \Col_Fill[6][5] ) );
  DLPQ3 \Col_Fill_reg[5][5]  ( .SN(n807), .D(n66440), .GN(n66380), .Q(
        \Col_Fill[5][5] ) );
  DLPQ3 \Col_Fill_reg[4][5]  ( .SN(n807), .D(n66440), .GN(n65560), .Q(
        \Col_Fill[4][5] ) );
  DLPQ3 \Col_Fill_reg[3][5]  ( .SN(n807), .D(n66440), .GN(n66378), .Q(
        \Col_Fill[3][5] ) );
  DLPQ3 \Col_Fill_reg[2][5]  ( .SN(n807), .D(n66440), .GN(n65558), .Q(
        \Col_Fill[2][5] ) );
  DLPQ3 \Col_Fill_reg[1][5]  ( .SN(n807), .D(n66440), .GN(n66376), .Q(
        \Col_Fill[1][5] ) );
  DLPQ3 \Col_Fill_reg[0][5]  ( .SN(n807), .D(n66440), .GN(n65556), .Q(
        \Col_Fill[0][5] ) );
  DLPQ3 \Col_Fill_reg[7][6]  ( .SN(n807), .D(n66441), .GN(n66382), .Q(
        \Col_Fill[7][6] ) );
  DLPQ3 \Col_Fill_reg[6][6]  ( .SN(n807), .D(n66441), .GN(n65562), .Q(
        \Col_Fill[6][6] ) );
  DLPQ3 \Col_Fill_reg[5][6]  ( .SN(n807), .D(n66441), .GN(n65561), .Q(
        \Col_Fill[5][6] ) );
  DLPQ3 \Col_Fill_reg[4][6]  ( .SN(n807), .D(n66441), .GN(n66379), .Q(
        \Col_Fill[4][6] ) );
  DLPQ3 \Col_Fill_reg[3][6]  ( .SN(n807), .D(n66441), .GN(n65559), .Q(
        \Col_Fill[3][6] ) );
  DLPQ3 \Col_Fill_reg[2][6]  ( .SN(n807), .D(n66441), .GN(n66377), .Q(
        \Col_Fill[2][6] ) );
  DLPQ3 \Col_Fill_reg[1][6]  ( .SN(n807), .D(n66441), .GN(n66376), .Q(
        \Col_Fill[1][6] ) );
  DLPQ3 \Col_Fill_reg[0][6]  ( .SN(n807), .D(n66441), .GN(n66375), .Q(
        \Col_Fill[0][6] ) );
  DLPQ3 \Col_Fill_reg[7][7]  ( .SN(n807), .D(n66442), .GN(n66382), .Q(
        \Col_Fill[7][7] ) );
  DLPQ3 \Col_Fill_reg[6][7]  ( .SN(n807), .D(n66442), .GN(n66381), .Q(
        \Col_Fill[6][7] ) );
  DLPQ3 \Col_Fill_reg[5][7]  ( .SN(n807), .D(n66442), .GN(n66380), .Q(
        \Col_Fill[5][7] ) );
  DLPQ3 \Col_Fill_reg[4][7]  ( .SN(n807), .D(n66442), .GN(n66379), .Q(
        \Col_Fill[4][7] ) );
  DLPQ3 \Col_Fill_reg[3][7]  ( .SN(n807), .D(n66442), .GN(n66378), .Q(
        \Col_Fill[3][7] ) );
  DLPQ3 \Col_Fill_reg[2][7]  ( .SN(n807), .D(n66442), .GN(n66377), .Q(
        \Col_Fill[2][7] ) );
  DLPQ3 \Col_Fill_reg[1][7]  ( .SN(n807), .D(n66442), .GN(n65557), .Q(
        \Col_Fill[1][7] ) );
  DLPQ3 \Col_Fill_reg[0][7]  ( .SN(n807), .D(n66442), .GN(n66375), .Q(
        \Col_Fill[0][7] ) );
  DLPQ3 \Col_Fill_reg[7][8]  ( .SN(n807), .D(n66443), .GN(n65563), .Q(
        \Col_Fill[7][8] ) );
  DLPQ3 \Col_Fill_reg[6][8]  ( .SN(n807), .D(n66443), .GN(n65562), .Q(
        \Col_Fill[6][8] ) );
  DLPQ3 \Col_Fill_reg[5][8]  ( .SN(n807), .D(n66443), .GN(n65561), .Q(
        \Col_Fill[5][8] ) );
  DLPQ3 \Col_Fill_reg[4][8]  ( .SN(n807), .D(n66443), .GN(n65560), .Q(
        \Col_Fill[4][8] ) );
  DLPQ3 \Col_Fill_reg[3][8]  ( .SN(n807), .D(n66443), .GN(n65559), .Q(
        \Col_Fill[3][8] ) );
  DLPQ3 \Col_Fill_reg[2][8]  ( .SN(n807), .D(n66443), .GN(n65558), .Q(
        \Col_Fill[2][8] ) );
  DLPQ3 \Col_Fill_reg[1][8]  ( .SN(n807), .D(n66443), .GN(n66376), .Q(
        \Col_Fill[1][8] ) );
  DLPQ3 \Col_Fill_reg[0][8]  ( .SN(n807), .D(n66443), .GN(n65556), .Q(
        \Col_Fill[0][8] ) );
  DLPQ3 \Col_Fill_reg[7][9]  ( .SN(n807), .D(n66444), .GN(n66382), .Q(
        \Col_Fill[7][9] ) );
  DLPQ3 \Col_Fill_reg[6][9]  ( .SN(n807), .D(n66444), .GN(n66381), .Q(
        \Col_Fill[6][9] ) );
  DLPQ3 \Col_Fill_reg[5][9]  ( .SN(n807), .D(n66444), .GN(n66380), .Q(
        \Col_Fill[5][9] ) );
  DLPQ3 \Col_Fill_reg[4][9]  ( .SN(n807), .D(n66444), .GN(n66379), .Q(
        \Col_Fill[4][9] ) );
  DLPQ3 \Col_Fill_reg[3][9]  ( .SN(n807), .D(n66444), .GN(n66378), .Q(
        \Col_Fill[3][9] ) );
  DLPQ3 \Col_Fill_reg[2][9]  ( .SN(n807), .D(n66444), .GN(n66377), .Q(
        \Col_Fill[2][9] ) );
  DLPQ3 \Col_Fill_reg[1][9]  ( .SN(n807), .D(n66444), .GN(n66376), .Q(
        \Col_Fill[1][9] ) );
  DLPQ3 \Col_Fill_reg[0][9]  ( .SN(n807), .D(n66444), .GN(n66375), .Q(
        \Col_Fill[0][9] ) );
  DLPQ3 \Col_Fill_reg[7][10]  ( .SN(n807), .D(n66445), .GN(n66382), .Q(
        \Col_Fill[7][10] ) );
  DLPQ3 \Col_Fill_reg[6][10]  ( .SN(n807), .D(n66445), .GN(n65562), .Q(
        \Col_Fill[6][10] ) );
  DLPQ3 \Col_Fill_reg[5][10]  ( .SN(n807), .D(n66445), .GN(n66380), .Q(
        \Col_Fill[5][10] ) );
  DLPQ3 \Col_Fill_reg[4][10]  ( .SN(n807), .D(n66445), .GN(n66379), .Q(
        \Col_Fill[4][10] ) );
  DLPQ3 \Col_Fill_reg[3][10]  ( .SN(n807), .D(n66445), .GN(n65559), .Q(
        \Col_Fill[3][10] ) );
  DLPQ3 \Col_Fill_reg[2][10]  ( .SN(n807), .D(n66445), .GN(n66377), .Q(
        \Col_Fill[2][10] ) );
  DLPQ3 \Col_Fill_reg[1][10]  ( .SN(n807), .D(n66445), .GN(n66376), .Q(
        \Col_Fill[1][10] ) );
  DLPQ3 \Col_Fill_reg[0][10]  ( .SN(n807), .D(n66445), .GN(n66375), .Q(
        \Col_Fill[0][10] ) );
  DLPQ3 \Col_Fill_reg[7][11]  ( .SN(n807), .D(n66446), .GN(n66382), .Q(
        \Col_Fill[7][11] ) );
  DLPQ3 \Col_Fill_reg[6][11]  ( .SN(n807), .D(n66446), .GN(n65562), .Q(
        \Col_Fill[6][11] ) );
  DLPQ3 \Col_Fill_reg[5][11]  ( .SN(n807), .D(n66446), .GN(n65561), .Q(
        \Col_Fill[5][11] ) );
  DLPQ3 \Col_Fill_reg[4][11]  ( .SN(n807), .D(n66446), .GN(n66379), .Q(
        \Col_Fill[4][11] ) );
  DLPQ3 \Col_Fill_reg[3][11]  ( .SN(n807), .D(n66446), .GN(n65559), .Q(
        \Col_Fill[3][11] ) );
  DLPQ3 \Col_Fill_reg[2][11]  ( .SN(n807), .D(n66446), .GN(n66377), .Q(
        \Col_Fill[2][11] ) );
  DLPQ3 \Col_Fill_reg[1][11]  ( .SN(n807), .D(n66446), .GN(n65557), .Q(
        \Col_Fill[1][11] ) );
  DLPQ3 \Col_Fill_reg[0][11]  ( .SN(n807), .D(n66446), .GN(n66375), .Q(
        \Col_Fill[0][11] ) );
  DLPQ3 \Col_Fill_reg[7][12]  ( .SN(n807), .D(n66447), .GN(n65563), .Q(
        \Col_Fill[7][12] ) );
  DLPQ3 \Col_Fill_reg[6][12]  ( .SN(n807), .D(n66447), .GN(n65562), .Q(
        \Col_Fill[6][12] ) );
  DLPQ3 \Col_Fill_reg[5][12]  ( .SN(n807), .D(n66447), .GN(n65561), .Q(
        \Col_Fill[5][12] ) );
  DLPQ3 \Col_Fill_reg[4][12]  ( .SN(n807), .D(n66447), .GN(n65560), .Q(
        \Col_Fill[4][12] ) );
  DLPQ3 \Col_Fill_reg[3][12]  ( .SN(n807), .D(n66447), .GN(n65559), .Q(
        \Col_Fill[3][12] ) );
  DLPQ3 \Col_Fill_reg[2][12]  ( .SN(n807), .D(n66447), .GN(n65558), .Q(
        \Col_Fill[2][12] ) );
  DLPQ3 \Col_Fill_reg[1][12]  ( .SN(n807), .D(n66447), .GN(n65557), .Q(
        \Col_Fill[1][12] ) );
  DLPQ3 \Col_Fill_reg[0][12]  ( .SN(n807), .D(n66447), .GN(n65556), .Q(
        \Col_Fill[0][12] ) );
  DLPQ3 \Col_Fill_reg[7][13]  ( .SN(n807), .D(n66448), .GN(n65563), .Q(
        \Col_Fill[7][13] ) );
  DLPQ3 \Col_Fill_reg[6][13]  ( .SN(n807), .D(n66448), .GN(n65562), .Q(
        \Col_Fill[6][13] ) );
  DLPQ3 \Col_Fill_reg[5][13]  ( .SN(n807), .D(n66448), .GN(n65561), .Q(
        \Col_Fill[5][13] ) );
  DLPQ3 \Col_Fill_reg[4][13]  ( .SN(n807), .D(n66448), .GN(n65560), .Q(
        \Col_Fill[4][13] ) );
  DLPQ3 \Col_Fill_reg[3][13]  ( .SN(n807), .D(n66448), .GN(n65559), .Q(
        \Col_Fill[3][13] ) );
  DLPQ3 \Col_Fill_reg[2][13]  ( .SN(n807), .D(n66448), .GN(n65558), .Q(
        \Col_Fill[2][13] ) );
  DLPQ3 \Col_Fill_reg[1][13]  ( .SN(n807), .D(n66448), .GN(n66376), .Q(
        \Col_Fill[1][13] ) );
  DLPQ3 \Col_Fill_reg[0][13]  ( .SN(n807), .D(n66448), .GN(n65556), .Q(
        \Col_Fill[0][13] ) );
  DLPQ3 \Col_Fill_reg[7][14]  ( .SN(n807), .D(n66449), .GN(n66382), .Q(
        \Col_Fill[7][14] ) );
  DLPQ3 \Col_Fill_reg[6][14]  ( .SN(n807), .D(n66449), .GN(n65562), .Q(
        \Col_Fill[6][14] ) );
  DLPQ3 \Col_Fill_reg[5][14]  ( .SN(n807), .D(n66449), .GN(n66380), .Q(
        \Col_Fill[5][14] ) );
  DLPQ3 \Col_Fill_reg[4][14]  ( .SN(n807), .D(n66449), .GN(n66379), .Q(
        \Col_Fill[4][14] ) );
  DLPQ3 \Col_Fill_reg[3][14]  ( .SN(n807), .D(n66449), .GN(n65559), .Q(
        \Col_Fill[3][14] ) );
  DLPQ3 \Col_Fill_reg[2][14]  ( .SN(n807), .D(n66449), .GN(n66377), .Q(
        \Col_Fill[2][14] ) );
  DLPQ3 \Col_Fill_reg[1][14]  ( .SN(n807), .D(n66449), .GN(n65557), .Q(
        \Col_Fill[1][14] ) );
  DLPQ3 \Col_Fill_reg[0][14]  ( .SN(n807), .D(n66449), .GN(n66375), .Q(
        \Col_Fill[0][14] ) );
  DLPQ3 \Col_Fill_reg[7][15]  ( .SN(n807), .D(n66450), .GN(n65563), .Q(
        \Col_Fill[7][15] ) );
  DLPQ3 \Col_Fill_reg[6][15]  ( .SN(n807), .D(n66450), .GN(n65562), .Q(
        \Col_Fill[6][15] ) );
  DLPQ3 \Col_Fill_reg[5][15]  ( .SN(n807), .D(n66450), .GN(n66380), .Q(
        \Col_Fill[5][15] ) );
  DLPQ3 \Col_Fill_reg[4][15]  ( .SN(n807), .D(n66450), .GN(n65560), .Q(
        \Col_Fill[4][15] ) );
  DLPQ3 \Col_Fill_reg[3][15]  ( .SN(n807), .D(n66450), .GN(n65559), .Q(
        \Col_Fill[3][15] ) );
  DLPQ3 \Col_Fill_reg[2][15]  ( .SN(n807), .D(n66450), .GN(n65558), .Q(
        \Col_Fill[2][15] ) );
  DLPQ3 \Col_Fill_reg[1][15]  ( .SN(n807), .D(n66450), .GN(n66376), .Q(
        \Col_Fill[1][15] ) );
  DLPQ3 \Col_Fill_reg[0][15]  ( .SN(n807), .D(n66450), .GN(n65556), .Q(
        \Col_Fill[0][15] ) );
  DLPQ3 \Col_Fill_reg[7][16]  ( .SN(n807), .D(n66451), .GN(n66382), .Q(
        \Col_Fill[7][16] ) );
  DLPQ3 \Col_Fill_reg[6][16]  ( .SN(n807), .D(n66451), .GN(n65562), .Q(
        \Col_Fill[6][16] ) );
  DLPQ3 \Col_Fill_reg[5][16]  ( .SN(n807), .D(n66451), .GN(n66380), .Q(
        \Col_Fill[5][16] ) );
  DLPQ3 \Col_Fill_reg[4][16]  ( .SN(n807), .D(n66451), .GN(n66379), .Q(
        \Col_Fill[4][16] ) );
  DLPQ3 \Col_Fill_reg[3][16]  ( .SN(n807), .D(n66451), .GN(n65559), .Q(
        \Col_Fill[3][16] ) );
  DLPQ3 \Col_Fill_reg[2][16]  ( .SN(n807), .D(n66451), .GN(n66377), .Q(
        \Col_Fill[2][16] ) );
  DLPQ3 \Col_Fill_reg[1][16]  ( .SN(n807), .D(n66451), .GN(n66376), .Q(
        \Col_Fill[1][16] ) );
  DLPQ3 \Col_Fill_reg[0][16]  ( .SN(n807), .D(n66451), .GN(n66375), .Q(
        \Col_Fill[0][16] ) );
  DLPQ3 \Col_Fill_reg[7][17]  ( .SN(n807), .D(n66452), .GN(n66382), .Q(
        \Col_Fill[7][17] ) );
  DLPQ3 \Col_Fill_reg[6][17]  ( .SN(n807), .D(n66452), .GN(n66381), .Q(
        \Col_Fill[6][17] ) );
  DLPQ3 \Col_Fill_reg[5][17]  ( .SN(n807), .D(n66452), .GN(n66380), .Q(
        \Col_Fill[5][17] ) );
  DLPQ3 \Col_Fill_reg[4][17]  ( .SN(n807), .D(n66452), .GN(n66379), .Q(
        \Col_Fill[4][17] ) );
  DLPQ3 \Col_Fill_reg[3][17]  ( .SN(n807), .D(n66452), .GN(n66378), .Q(
        \Col_Fill[3][17] ) );
  DLPQ3 \Col_Fill_reg[2][17]  ( .SN(n807), .D(n66452), .GN(n66377), .Q(
        \Col_Fill[2][17] ) );
  DLPQ3 \Col_Fill_reg[1][17]  ( .SN(n807), .D(n66452), .GN(n65557), .Q(
        \Col_Fill[1][17] ) );
  DLPQ3 \Col_Fill_reg[0][17]  ( .SN(n807), .D(n66452), .GN(n66375), .Q(
        \Col_Fill[0][17] ) );
  DLPQ3 \Col_Fill_reg[7][18]  ( .SN(n807), .D(n66453), .GN(n65563), .Q(
        \Col_Fill[7][18] ) );
  DLPQ3 \Col_Fill_reg[6][18]  ( .SN(n807), .D(n66453), .GN(n66381), .Q(
        \Col_Fill[6][18] ) );
  DLPQ3 \Col_Fill_reg[5][18]  ( .SN(n807), .D(n66453), .GN(n65561), .Q(
        \Col_Fill[5][18] ) );
  DLPQ3 \Col_Fill_reg[4][18]  ( .SN(n807), .D(n66453), .GN(n65560), .Q(
        \Col_Fill[4][18] ) );
  DLPQ3 \Col_Fill_reg[3][18]  ( .SN(n807), .D(n66453), .GN(n66378), .Q(
        \Col_Fill[3][18] ) );
  DLPQ3 \Col_Fill_reg[2][18]  ( .SN(n807), .D(n66453), .GN(n65558), .Q(
        \Col_Fill[2][18] ) );
  DLPQ3 \Col_Fill_reg[1][18]  ( .SN(n807), .D(n66453), .GN(n66376), .Q(
        \Col_Fill[1][18] ) );
  DLPQ3 \Col_Fill_reg[0][18]  ( .SN(n807), .D(n66453), .GN(n65556), .Q(
        \Col_Fill[0][18] ) );
  DLPQ3 \Col_Fill_reg[7][19]  ( .SN(n807), .D(n66454), .GN(n66382), .Q(
        \Col_Fill[7][19] ) );
  DLPQ3 \Col_Fill_reg[6][19]  ( .SN(n807), .D(n66454), .GN(n66381), .Q(
        \Col_Fill[6][19] ) );
  DLPQ3 \Col_Fill_reg[5][19]  ( .SN(n807), .D(n66454), .GN(n66380), .Q(
        \Col_Fill[5][19] ) );
  DLPQ3 \Col_Fill_reg[4][19]  ( .SN(n807), .D(n66454), .GN(n66379), .Q(
        \Col_Fill[4][19] ) );
  DLPQ3 \Col_Fill_reg[3][19]  ( .SN(n807), .D(n66454), .GN(n66378), .Q(
        \Col_Fill[3][19] ) );
  DLPQ3 \Col_Fill_reg[2][19]  ( .SN(n807), .D(n66454), .GN(n66377), .Q(
        \Col_Fill[2][19] ) );
  DLPQ3 \Col_Fill_reg[1][19]  ( .SN(n807), .D(n66454), .GN(n65557), .Q(
        \Col_Fill[1][19] ) );
  DLPQ3 \Col_Fill_reg[0][19]  ( .SN(n807), .D(n66454), .GN(n66375), .Q(
        \Col_Fill[0][19] ) );
  DLPQ3 \Col_Fill_reg[7][20]  ( .SN(n807), .D(n66455), .GN(n65563), .Q(
        \Col_Fill[7][20] ) );
  DLPQ3 \Col_Fill_reg[6][20]  ( .SN(n807), .D(n66455), .GN(n65562), .Q(
        \Col_Fill[6][20] ) );
  DLPQ3 \Col_Fill_reg[5][20]  ( .SN(n807), .D(n66455), .GN(n65561), .Q(
        \Col_Fill[5][20] ) );
  DLPQ3 \Col_Fill_reg[4][20]  ( .SN(n807), .D(n66455), .GN(n65560), .Q(
        \Col_Fill[4][20] ) );
  DLPQ3 \Col_Fill_reg[3][20]  ( .SN(n807), .D(n66455), .GN(n65559), .Q(
        \Col_Fill[3][20] ) );
  DLPQ3 \Col_Fill_reg[2][20]  ( .SN(n807), .D(n66455), .GN(n65558), .Q(
        \Col_Fill[2][20] ) );
  DLPQ3 \Col_Fill_reg[1][20]  ( .SN(n807), .D(n66455), .GN(n66376), .Q(
        \Col_Fill[1][20] ) );
  DLPQ3 \Col_Fill_reg[0][20]  ( .SN(n807), .D(n66455), .GN(n65556), .Q(
        \Col_Fill[0][20] ) );
  DLPQ3 \Col_Fill_reg[7][21]  ( .SN(n807), .D(n66456), .GN(n66382), .Q(
        \Col_Fill[7][21] ) );
  DLPQ3 \Col_Fill_reg[6][21]  ( .SN(n807), .D(n66456), .GN(n66381), .Q(
        \Col_Fill[6][21] ) );
  DLPQ3 \Col_Fill_reg[5][21]  ( .SN(n807), .D(n66456), .GN(n65561), .Q(
        \Col_Fill[5][21] ) );
  DLPQ3 \Col_Fill_reg[4][21]  ( .SN(n807), .D(n66456), .GN(n66379), .Q(
        \Col_Fill[4][21] ) );
  DLPQ3 \Col_Fill_reg[3][21]  ( .SN(n807), .D(n66456), .GN(n66378), .Q(
        \Col_Fill[3][21] ) );
  DLPQ3 \Col_Fill_reg[2][21]  ( .SN(n807), .D(n66456), .GN(n66377), .Q(
        \Col_Fill[2][21] ) );
  DLPQ3 \Col_Fill_reg[1][21]  ( .SN(n807), .D(n66456), .GN(n65557), .Q(
        \Col_Fill[1][21] ) );
  DLPQ3 \Col_Fill_reg[0][21]  ( .SN(n807), .D(n66456), .GN(n66375), .Q(
        \Col_Fill[0][21] ) );
  DLPQ3 \Col_Fill_reg[7][22]  ( .SN(n807), .D(n66457), .GN(n65563), .Q(
        \Col_Fill[7][22] ) );
  DLPQ3 \Col_Fill_reg[6][22]  ( .SN(n807), .D(n66457), .GN(n65562), .Q(
        \Col_Fill[6][22] ) );
  DLPQ3 \Col_Fill_reg[5][22]  ( .SN(n807), .D(n66457), .GN(n66380), .Q(
        \Col_Fill[5][22] ) );
  DLPQ3 \Col_Fill_reg[4][22]  ( .SN(n807), .D(n66457), .GN(n65560), .Q(
        \Col_Fill[4][22] ) );
  DLPQ3 \Col_Fill_reg[3][22]  ( .SN(n807), .D(n66457), .GN(n65559), .Q(
        \Col_Fill[3][22] ) );
  DLPQ3 \Col_Fill_reg[2][22]  ( .SN(n807), .D(n66457), .GN(n65558), .Q(
        \Col_Fill[2][22] ) );
  DLPQ3 \Col_Fill_reg[1][22]  ( .SN(n807), .D(n66457), .GN(n66376), .Q(
        \Col_Fill[1][22] ) );
  DLPQ3 \Col_Fill_reg[0][22]  ( .SN(n807), .D(n66457), .GN(n65556), .Q(
        \Col_Fill[0][22] ) );
  DLPQ3 \Col_Fill_reg[7][23]  ( .SN(n807), .D(n66458), .GN(n66382), .Q(
        \Col_Fill[7][23] ) );
  DLPQ3 \Col_Fill_reg[6][23]  ( .SN(n807), .D(n66458), .GN(n66381), .Q(
        \Col_Fill[6][23] ) );
  DLPQ3 \Col_Fill_reg[5][23]  ( .SN(n807), .D(n66458), .GN(n66380), .Q(
        \Col_Fill[5][23] ) );
  DLPQ3 \Col_Fill_reg[4][23]  ( .SN(n807), .D(n66458), .GN(n66379), .Q(
        \Col_Fill[4][23] ) );
  DLPQ3 \Col_Fill_reg[3][23]  ( .SN(n807), .D(n66458), .GN(n66378), .Q(
        \Col_Fill[3][23] ) );
  DLPQ3 \Col_Fill_reg[2][23]  ( .SN(n807), .D(n66458), .GN(n66377), .Q(
        \Col_Fill[2][23] ) );
  DLPQ3 \Col_Fill_reg[1][23]  ( .SN(n807), .D(n66458), .GN(n65557), .Q(
        \Col_Fill[1][23] ) );
  DLPQ3 \Col_Fill_reg[0][23]  ( .SN(n807), .D(n66458), .GN(n66375), .Q(
        \Col_Fill[0][23] ) );
  DLPQ3 \Col_Fill_reg[7][24]  ( .SN(n807), .D(n66459), .GN(n65563), .Q(
        \Col_Fill[7][24] ) );
  DLPQ3 \Col_Fill_reg[6][24]  ( .SN(n807), .D(n66459), .GN(n66381), .Q(
        \Col_Fill[6][24] ) );
  DLPQ3 \Col_Fill_reg[5][24]  ( .SN(n807), .D(n66459), .GN(n66380), .Q(
        \Col_Fill[5][24] ) );
  DLPQ3 \Col_Fill_reg[4][24]  ( .SN(n807), .D(n66459), .GN(n65560), .Q(
        \Col_Fill[4][24] ) );
  DLPQ3 \Col_Fill_reg[3][24]  ( .SN(n807), .D(n66459), .GN(n66378), .Q(
        \Col_Fill[3][24] ) );
  DLPQ3 \Col_Fill_reg[2][24]  ( .SN(n807), .D(n66459), .GN(n65558), .Q(
        \Col_Fill[2][24] ) );
  DLPQ3 \Col_Fill_reg[1][24]  ( .SN(n807), .D(n66459), .GN(n65557), .Q(
        \Col_Fill[1][24] ) );
  DLPQ3 \Col_Fill_reg[0][24]  ( .SN(n807), .D(n66459), .GN(n65556), .Q(
        \Col_Fill[0][24] ) );
  DLPQ3 \Col_Fill_reg[7][25]  ( .SN(n807), .D(n66460), .GN(n65563), .Q(
        \Col_Fill[7][25] ) );
  DLPQ3 \Col_Fill_reg[6][25]  ( .SN(n807), .D(n66460), .GN(n65562), .Q(
        \Col_Fill[6][25] ) );
  DLPQ3 \Col_Fill_reg[5][25]  ( .SN(n807), .D(n66460), .GN(n65561), .Q(
        \Col_Fill[5][25] ) );
  DLPQ3 \Col_Fill_reg[4][25]  ( .SN(n807), .D(n66460), .GN(n65560), .Q(
        \Col_Fill[4][25] ) );
  DLPQ3 \Col_Fill_reg[3][25]  ( .SN(n807), .D(n66460), .GN(n65559), .Q(
        \Col_Fill[3][25] ) );
  DLPQ3 \Col_Fill_reg[2][25]  ( .SN(n807), .D(n66460), .GN(n65558), .Q(
        \Col_Fill[2][25] ) );
  DLPQ3 \Col_Fill_reg[1][25]  ( .SN(n807), .D(n66460), .GN(n65557), .Q(
        \Col_Fill[1][25] ) );
  DLPQ3 \Col_Fill_reg[0][25]  ( .SN(n807), .D(n66460), .GN(n65556), .Q(
        \Col_Fill[0][25] ) );
  DLPQ3 \Col_Fill_reg[7][26]  ( .SN(n807), .D(n66461), .GN(n65563), .Q(
        \Col_Fill[7][26] ) );
  DLPQ3 \Col_Fill_reg[6][26]  ( .SN(n807), .D(n66461), .GN(n66381), .Q(
        \Col_Fill[6][26] ) );
  DLPQ3 \Col_Fill_reg[5][26]  ( .SN(n807), .D(n66461), .GN(n66380), .Q(
        \Col_Fill[5][26] ) );
  DLPQ3 \Col_Fill_reg[4][26]  ( .SN(n807), .D(n66461), .GN(n65560), .Q(
        \Col_Fill[4][26] ) );
  DLPQ3 \Col_Fill_reg[3][26]  ( .SN(n807), .D(n66461), .GN(n66378), .Q(
        \Col_Fill[3][26] ) );
  DLPQ3 \Col_Fill_reg[2][26]  ( .SN(n807), .D(n66461), .GN(n65558), .Q(
        \Col_Fill[2][26] ) );
  DLPQ3 \Col_Fill_reg[1][26]  ( .SN(n807), .D(n66461), .GN(n65557), .Q(
        \Col_Fill[1][26] ) );
  DLPQ3 \Col_Fill_reg[0][26]  ( .SN(n807), .D(n66461), .GN(n65556), .Q(
        \Col_Fill[0][26] ) );
  DLPQ3 \Col_Fill_reg[7][27]  ( .SN(n807), .D(n66462), .GN(n65563), .Q(
        \Col_Fill[7][27] ) );
  DLPQ3 \Col_Fill_reg[6][27]  ( .SN(n807), .D(n66462), .GN(n66381), .Q(
        \Col_Fill[6][27] ) );
  DLPQ3 \Col_Fill_reg[5][27]  ( .SN(n807), .D(n66462), .GN(n65561), .Q(
        \Col_Fill[5][27] ) );
  DLPQ3 \Col_Fill_reg[4][27]  ( .SN(n807), .D(n66462), .GN(n65560), .Q(
        \Col_Fill[4][27] ) );
  DLPQ3 \Col_Fill_reg[3][27]  ( .SN(n807), .D(n66462), .GN(n66378), .Q(
        \Col_Fill[3][27] ) );
  DLPQ3 \Col_Fill_reg[2][27]  ( .SN(n807), .D(n66462), .GN(n65558), .Q(
        \Col_Fill[2][27] ) );
  DLPQ3 \Col_Fill_reg[1][27]  ( .SN(n807), .D(n66462), .GN(n65557), .Q(
        \Col_Fill[1][27] ) );
  DLPQ3 \Col_Fill_reg[0][27]  ( .SN(n807), .D(n66462), .GN(n65556), .Q(
        \Col_Fill[0][27] ) );
  DLPQ3 \Col_Fill_reg[7][28]  ( .SN(n807), .D(n66463), .GN(n65563), .Q(
        \Col_Fill[7][28] ) );
  DLPQ3 \Col_Fill_reg[6][28]  ( .SN(n807), .D(n66463), .GN(n66381), .Q(
        \Col_Fill[6][28] ) );
  DLPQ3 \Col_Fill_reg[5][28]  ( .SN(n807), .D(n66463), .GN(n66380), .Q(
        \Col_Fill[5][28] ) );
  DLPQ3 \Col_Fill_reg[4][28]  ( .SN(n807), .D(n66463), .GN(n65560), .Q(
        \Col_Fill[4][28] ) );
  DLPQ3 \Col_Fill_reg[3][28]  ( .SN(n807), .D(n66463), .GN(n66378), .Q(
        \Col_Fill[3][28] ) );
  DLPQ3 \Col_Fill_reg[2][28]  ( .SN(n807), .D(n66463), .GN(n65558), .Q(
        \Col_Fill[2][28] ) );
  DLPQ3 \Col_Fill_reg[1][28]  ( .SN(n807), .D(n66463), .GN(n65557), .Q(
        \Col_Fill[1][28] ) );
  DLPQ3 \Col_Fill_reg[0][28]  ( .SN(n807), .D(n66463), .GN(n65556), .Q(
        \Col_Fill[0][28] ) );
  DLPQ3 \Col_Fill_reg[7][29]  ( .SN(n807), .D(n66464), .GN(n65563), .Q(
        \Col_Fill[7][29] ) );
  DLPQ3 \Col_Fill_reg[6][29]  ( .SN(n807), .D(n66464), .GN(n65562), .Q(
        \Col_Fill[6][29] ) );
  DLPQ3 \Col_Fill_reg[5][29]  ( .SN(n807), .D(n66464), .GN(n65561), .Q(
        \Col_Fill[5][29] ) );
  DLPQ3 \Col_Fill_reg[4][29]  ( .SN(n807), .D(n66464), .GN(n65560), .Q(
        \Col_Fill[4][29] ) );
  DLPQ3 \Col_Fill_reg[3][29]  ( .SN(n807), .D(n66464), .GN(n65559), .Q(
        \Col_Fill[3][29] ) );
  DLPQ3 \Col_Fill_reg[2][29]  ( .SN(n807), .D(n66464), .GN(n65558), .Q(
        \Col_Fill[2][29] ) );
  DLPQ3 \Col_Fill_reg[1][29]  ( .SN(n807), .D(n66464), .GN(n65557), .Q(
        \Col_Fill[1][29] ) );
  DLPQ3 \Col_Fill_reg[0][29]  ( .SN(n807), .D(n66464), .GN(n65556), .Q(
        \Col_Fill[0][29] ) );
  DLPQ3 \Col_Fill_reg[7][30]  ( .SN(n807), .D(n66465), .GN(n65563), .Q(
        \Col_Fill[7][30] ) );
  DLPQ3 \Col_Fill_reg[6][30]  ( .SN(n807), .D(n66465), .GN(n65562), .Q(
        \Col_Fill[6][30] ) );
  DLPQ3 \Col_Fill_reg[5][30]  ( .SN(n807), .D(n66465), .GN(n66380), .Q(
        \Col_Fill[5][30] ) );
  DLPQ3 \Col_Fill_reg[4][30]  ( .SN(n807), .D(n66465), .GN(n65560), .Q(
        \Col_Fill[4][30] ) );
  DLPQ3 \Col_Fill_reg[3][30]  ( .SN(n807), .D(n66465), .GN(n65559), .Q(
        \Col_Fill[3][30] ) );
  DLPQ3 \Col_Fill_reg[2][30]  ( .SN(n807), .D(n66465), .GN(n65558), .Q(
        \Col_Fill[2][30] ) );
  DLPQ3 \Col_Fill_reg[0][30]  ( .SN(n807), .D(n66465), .GN(n65556), .Q(
        \Col_Fill[0][30] ) );
  DLPQ3 \n_reg[0]  ( .SN(n807), .D(n66431), .GN(n65564), .Q(N1207) );
  DLPQ3 \n_reg[1]  ( .SN(n807), .D(n66430), .GN(n65564), .Q(N1208) );
  DLPQ3 \n_reg[2]  ( .SN(n807), .D(n66429), .GN(n65564), .Q(N1167) );
  DLPQ3 \n_reg[3]  ( .SN(n807), .D(n66428), .GN(n66393), .Q(n[3]) );
  DLPQ3 \n_reg[4]  ( .SN(n807), .D(n66427), .GN(n66393), .Q(n[4]) );
  DLPQ3 \n_reg[5]  ( .SN(n807), .D(n66426), .GN(n66393), .Q(n[5]) );
  DLPQ3 \n_reg[6]  ( .SN(n807), .D(n66425), .GN(n65564), .Q(n[6]) );
  DLPQ3 \n_reg[7]  ( .SN(n807), .D(n66424), .GN(n66393), .Q(n[7]) );
  DLPQ3 \n_reg[8]  ( .SN(n807), .D(n66423), .GN(n66393), .Q(n[8]) );
  DLPQ3 \n_reg[9]  ( .SN(n807), .D(n66422), .GN(n66393), .Q(n[9]) );
  DLPQ3 \n_reg[10]  ( .SN(n807), .D(n66421), .GN(n65564), .Q(n[10]) );
  DLPQ3 \n_reg[11]  ( .SN(n807), .D(n66420), .GN(n66393), .Q(n[11]) );
  DLPQ3 \n_reg[12]  ( .SN(n807), .D(n66419), .GN(n66393), .Q(n[12]) );
  DLPQ3 \n_reg[13]  ( .SN(n807), .D(n66418), .GN(n65564), .Q(n[13]) );
  DLPQ3 \n_reg[14]  ( .SN(n807), .D(n66417), .GN(n66393), .Q(n[14]) );
  DLPQ3 \n_reg[15]  ( .SN(n807), .D(n66416), .GN(n66393), .Q(n[15]) );
  DLPQ3 \n_reg[16]  ( .SN(n807), .D(n66415), .GN(n65564), .Q(n[16]) );
  DLPQ3 \n_reg[17]  ( .SN(n807), .D(n66414), .GN(n65564), .Q(n[17]) );
  DLPQ3 \n_reg[18]  ( .SN(n807), .D(n66413), .GN(n66393), .Q(n[18]) );
  DLPQ3 \n_reg[19]  ( .SN(n807), .D(n66412), .GN(n66393), .Q(n[19]) );
  DLPQ3 \n_reg[20]  ( .SN(n807), .D(n66411), .GN(n65564), .Q(n[20]) );
  DLPQ3 \n_reg[21]  ( .SN(n807), .D(n66410), .GN(n66393), .Q(n[21]) );
  DLPQ3 \n_reg[22]  ( .SN(n807), .D(n66409), .GN(n65564), .Q(n[22]) );
  DLPQ3 \n_reg[23]  ( .SN(n807), .D(n66408), .GN(n66393), .Q(n[23]) );
  DLPQ3 \n_reg[24]  ( .SN(n807), .D(n66407), .GN(n65564), .Q(n[24]) );
  DLPQ3 \n_reg[25]  ( .SN(n807), .D(n66406), .GN(n65564), .Q(n[25]) );
  DLPQ3 \n_reg[26]  ( .SN(n807), .D(n66405), .GN(n65564), .Q(n[26]) );
  DLPQ3 \n_reg[27]  ( .SN(n807), .D(n66404), .GN(n65564), .Q(n[27]) );
  DLPQ3 \n_reg[28]  ( .SN(n807), .D(n66403), .GN(n65564), .Q(n[28]) );
  DLPQ3 \n_reg[29]  ( .SN(n807), .D(n66402), .GN(n65564), .Q(n[29]) );
  DLPQ3 \n_reg[30]  ( .SN(n807), .D(n66401), .GN(n65564), .Q(n[30]) );
  DLPQ3 \n_reg[31]  ( .SN(n807), .D(n66400), .GN(n65564), .Q(n[31]) );
  DF3 \C4_OUT_reg[1]  ( .D(n65434), .C(CLK), .Q(C4_OUT[1]), .QN(n1681) );
  DLPQ3 \LED_PIN_reg[22]  ( .SN(n807), .D(N2677), .GN(n66360), .Q(LED_PIN[22])
         );
  DLPQ3 \LED_PIN_reg[11]  ( .SN(n807), .D(N2655), .GN(n66344), .Q(LED_PIN[11])
         );
  DLPQ3 \LED_PIN_reg[8]  ( .SN(n807), .D(N2649), .GN(n66341), .Q(LED_PIN[8])
         );
  DLPQ3 \LED_PIN_reg[5]  ( .SN(n807), .D(N2643), .GN(n66350), .Q(LED_PIN[5])
         );
  DLPQ3 \LED_PIN_reg[2]  ( .SN(n807), .D(N2637), .GN(n66337), .Q(LED_PIN[2])
         );
  DLPQ3 \LED_PIN_reg[19]  ( .SN(n807), .D(N2671), .GN(n66348), .Q(LED_PIN[19])
         );
  DLPQ3 \LED_PIN_reg[16]  ( .SN(n807), .D(N2665), .GN(n66345), .Q(LED_PIN[16])
         );
  DLPQ3 \LED_PIN_reg[13]  ( .SN(n807), .D(N2659), .GN(n66355), .Q(LED_PIN[13])
         );
  DLPQ3 \LED_PIN_reg[10]  ( .SN(n807), .D(N2653), .GN(n66343), .Q(LED_PIN[10])
         );
  DLPQ3 \LED_PIN_reg[7]  ( .SN(n807), .D(N2647), .GN(n66353), .Q(LED_PIN[7])
         );
  DLPQ3 \LED_PIN_reg[4]  ( .SN(n807), .D(N2641), .GN(n66349), .Q(LED_PIN[4])
         );
  DLPQ3 \LED_PIN_reg[1]  ( .SN(n807), .D(N2635), .GN(n66336), .Q(LED_PIN[1])
         );
  DLPQ3 \LED_PIN_reg[23]  ( .SN(n807), .D(N2679), .GN(n66361), .Q(LED_PIN[23])
         );
  DLPQ3 \LED_PIN_reg[20]  ( .SN(n807), .D(N2673), .GN(n66358), .Q(LED_PIN[20])
         );
  DLPQ3 \LED_PIN_reg[17]  ( .SN(n807), .D(N2667), .GN(n66346), .Q(LED_PIN[17])
         );
  DLPQ3 \LED_PIN_reg[14]  ( .SN(n807), .D(N2661), .GN(n66356), .Q(LED_PIN[14])
         );
  DLPQ3 \LED_PIN_reg[21]  ( .SN(n807), .D(N2675), .GN(n66359), .Q(LED_PIN[21])
         );
  DLPQ3 \LED_PIN_reg[18]  ( .SN(n807), .D(N2669), .GN(n66347), .Q(LED_PIN[18])
         );
  DLPQ3 \LED_PIN_reg[15]  ( .SN(n807), .D(N2663), .GN(n66357), .Q(LED_PIN[15])
         );
  DLPQ3 \LED_PIN_reg[12]  ( .SN(n807), .D(N2657), .GN(n66354), .Q(LED_PIN[12])
         );
  DLPQ3 \LED_PIN_reg[9]  ( .SN(n807), .D(N2651), .GN(n66342), .Q(LED_PIN[9])
         );
  DLPQ3 \LED_PIN_reg[6]  ( .SN(n807), .D(N2645), .GN(n66352), .Q(LED_PIN[6])
         );
  DLPQ3 \LED_PIN_reg[3]  ( .SN(n807), .D(N2639), .GN(n66339), .Q(LED_PIN[3])
         );
  DLPQ3 \LED_PIN_reg[0]  ( .SN(n807), .D(N2633), .GN(n66334), .Q(LED_PIN[0])
         );
  Connect4_DW01_add_97 add_0_root_sub_0_root_sub_136_2 ( .A({n65541, n65540, 
        n65540, n65540, n65540, n65541, n65541, n65541, n65541, n65540, n65540, 
        n65540, n65540, n65541, n65541, n65541, n65541, n65540, n65540, n65540, 
        n65540, n65541, n65541, N1380, N1379, N1378, N1377, N1376, n65741, 
        n807, n807, n807}), .B({N1331, N1330, N1329, N1328, N1327, N1326, 
        N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, 
        N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, 
        N1305, N1304, N1303, N1302, N1301, n65546}), .CI(n65544), .SUM({N1435, 
        N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, 
        N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, 
        N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, 
        N1404}) );
  Connect4_DW01_add_96 add_0_root_sub_0_root_sub_167_2 ( .A({n65543, N1946, 
        n65543, N1946, n65543, n65543, n65543, n65543, n65543, N1946, n65543, 
        N1946, n65543, n65543, n65543, n65543, n65543, n65543, n65543, n65543, 
        n65543, n65543, n65543, N1923, N1922, N1921, N1920, N1919, n65740, 
        n807, n807, n807}), .B({N1874, N1873, N1872, N1871, N1870, N1869, 
        N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, 
        N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, 
        N1848, N1847, N1846, N1845, N1844, n65545}), .CI(n65544), .SUM({N1978, 
        N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, 
        N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, 
        N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, 
        N1947}) );
  ADD22 \add_1_root_add_157_3/U1_1_1  ( .A(O_play[1]), .B(n65419), .CO(
        \add_1_root_add_157_3/carry[2] ), .S(N1836) );
  ADD22 \add_1_root_add_157_3/U1_1_2  ( .A(O_play[2]), .B(
        \add_1_root_add_157_3/carry[2] ), .CO(N1838), .S(N1837) );
  ADD32 \add_0_root_sub_0_root_sub_297_3/U1_3  ( .A(n65593), .B(n65581), .CI(
        \add_0_root_sub_0_root_sub_297_3/carry [3]), .CO(
        \add_0_root_sub_0_root_sub_297_3/carry [4]), .S(N694) );
  ADD32 \add_0_root_sub_0_root_sub_297_3/U1_4  ( .A(n65597), .B(N2901), .CI(
        \add_0_root_sub_0_root_sub_297_3/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_297_3/carry [5]), .S(N695) );
  ADD32 \add_0_root_sub_0_root_sub_297_6/U1_3  ( .A(n65593), .B(n65579), .CI(
        \add_0_root_sub_0_root_sub_297_6/carry [3]), .CO(
        \add_0_root_sub_0_root_sub_297_6/carry [4]), .S(N700) );
  ADD32 \add_0_root_sub_0_root_sub_297_6/U1_4  ( .A(n65597), .B(N2919), .CI(
        \add_0_root_sub_0_root_sub_297_6/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_297_6/carry [5]), .S(N701) );
  ADD32 \add_0_root_sub_0_root_sub_297_9/U1_4  ( .A(m[1]), .B(N2937), .CI(
        \add_0_root_sub_0_root_sub_297_9/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_297_9/carry [5]), .S(N707) );
  ADD32 \add_0_root_sub_0_root_sub_369_3/U1_4  ( .A(n65605), .B(N5171), .CI(
        \add_0_root_sub_0_root_sub_369_3/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_369_3/carry [5]), .S(N983) );
  ADD32 \add_0_root_sub_0_root_sub_369_6/U1_4  ( .A(N5183), .B(N5189), .CI(
        \add_0_root_sub_0_root_sub_369_6/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_369_6/carry [5]), .S(N989) );
  ADD32 \add_0_root_sub_0_root_sub_369_9/U1_4  ( .A(m[1]), .B(N5207), .CI(
        \add_0_root_sub_0_root_sub_369_9/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_369_9/carry [5]), .S(N995) );
  ADD32 \add_0_root_sub_0_root_sub_300_5/U1_4  ( .A(n65605), .B(N3073), .CI(
        \add_0_root_sub_0_root_sub_300_5/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_300_5/carry [5]), .S(N719) );
  ADD32 \add_0_root_sub_0_root_sub_300_8/U1_4  ( .A(N3085), .B(N3091), .CI(
        \add_0_root_sub_0_root_sub_300_8/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_300_8/carry [5]), .S(N725) );
  ADD32 \add_0_root_sub_0_root_sub_372_5/U1_4  ( .A(n65605), .B(N5343), .CI(
        \add_0_root_sub_0_root_sub_372_5/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_372_5/carry [5]), .S(N1007) );
  ADD32 \add_0_root_sub_0_root_sub_372_8/U1_4  ( .A(N5355), .B(N5361), .CI(
        \add_0_root_sub_0_root_sub_372_8/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_372_8/carry [5]), .S(N1013) );
  ADD32 \add_0_root_sub_0_root_sub_303_7/U1_4  ( .A(n65605), .B(N3246), .CI(
        \add_0_root_sub_0_root_sub_303_7/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_303_7/carry [5]), .S(N743) );
  ADD32 \add_0_root_sub_0_root_sub_375_7/U1_4  ( .A(n65608), .B(N5516), .CI(
        \add_0_root_sub_0_root_sub_375_7/carry [4]), .CO(
        \add_0_root_sub_0_root_sub_375_7/carry [5]), .S(N1031) );
  ADD32 \r11558/U1_4  ( .A(N3510), .B(N11267), .CI(\r11558/carry [4]), .CO(
        \r11558/carry [5]), .S(N1067) );
  ADD32 \r11557/U1_4  ( .A(N3510), .B(N11261), .CI(\r11557/carry [4]), .CO(
        \r11557/carry [5]), .S(N1061) );
  ADD32 \r11556/U1_4  ( .A(N3510), .B(N11255), .CI(\r11556/carry [4]), .CO(
        \r11556/carry [5]), .S(N1055) );
  ADD32 \r12191/U1_4  ( .A(N3637), .B(N11291), .CI(\r12191/carry [4]), .CO(
        \r12191/carry [5]), .S(N1085) );
  ADD32 \r12190/U1_4  ( .A(N3637), .B(N11285), .CI(\r12190/carry [4]), .CO(
        \r12190/carry [5]), .S(N1079) );
  ADD32 \r12187/U1_4  ( .A(N3637), .B(n65597), .CI(\r32996/carry [4]), .CO(
        \r12187/carry[5] ), .S(N1073) );
  ADD22 \r13451/U1_1_1  ( .A(n65757), .B(n65839), .CO(\r13451/carry [2]), .S(
        N1112) );
  ADD22 \r13451/U1_1_2  ( .A(n65918), .B(\r13451/carry [2]), .CO(
        \r13451/carry [3]), .S(N1113) );
  ADD22 \r13451/U1_1_3  ( .A(N11412), .B(\r13451/carry [3]), .CO(
        \r13451/carry [4]), .S(N1114) );
  ADD22 \r13451/U1_1_4  ( .A(N1121), .B(\r13451/carry [4]), .CO(
        \r13451/carry [5]), .S(N1115) );
  ADD32 \r13450/U1_4  ( .A(N3899), .B(N11321), .CI(\r13450/carry [4]), .CO(
        \r13450/carry [5]), .S(N1109) );
  ADD32 \r13449/U1_4  ( .A(N3899), .B(n65597), .CI(\r32996/carry [4]), .CO(
        \r13449/carry[5] ), .S(N1121) );
  ADD32 \add_0_root_add_0_root_sub_325_4_cf/U1_3  ( .A(n65593), .B(n65585), 
        .CI(\add_0_root_add_0_root_sub_325_4_cf/carry [3]), .CO(
        \add_0_root_add_0_root_sub_325_4_cf/carry [4]), .S(N838) );
  ADD32 \add_0_root_add_0_root_sub_325_4_cf/U1_4  ( .A(n65597), .B(N11351), 
        .CI(\add_0_root_add_0_root_sub_325_4_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_325_4_cf/carry [5]), .S(N839) );
  ADD32 \add_0_root_add_0_root_sub_325_8_cf/U1_3  ( .A(n65593), .B(N3200), 
        .CI(\add_0_root_add_0_root_sub_325_8_cf/carry [3]), .CO(
        \add_0_root_add_0_root_sub_325_8_cf/carry [4]), .S(N844) );
  ADD32 \add_0_root_add_0_root_sub_325_8_cf/U1_4  ( .A(n65597), .B(N11357), 
        .CI(\add_0_root_add_0_root_sub_325_8_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_325_8_cf/carry [5]), .S(N845) );
  ADD32 \add_0_root_add_0_root_sub_325_12_cf/U1_3  ( .A(n65593), .B(n65584), 
        .CI(n65915), .CO(\add_0_root_add_0_root_sub_325_12_cf/carry [4]), .S(
        N850) );
  ADD32 \add_0_root_add_0_root_sub_325_12_cf/U1_4  ( .A(n65597), .B(N11363), 
        .CI(\add_0_root_add_0_root_sub_325_12_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_325_12_cf/carry [5]), .S(N851) );
  ADD32 \add_0_root_add_0_root_sub_397_4_cf/U1_4  ( .A(n65608), .B(N11333), 
        .CI(\add_0_root_add_0_root_sub_397_4_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_397_4_cf/carry [5]), .S(N1127) );
  ADD32 \add_0_root_add_0_root_sub_397_8_cf/U1_4  ( .A(N6311), .B(N11339), 
        .CI(\add_0_root_add_0_root_sub_397_8_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_397_8_cf/carry [5]), .S(N1133) );
  ADD32 \add_0_root_add_0_root_sub_397_12_cf/U1_4  ( .A(m[1]), .B(N11345), 
        .CI(\add_0_root_add_0_root_sub_397_12_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_397_12_cf/carry [5]), .S(N1139) );
  ADD32 \add_0_root_add_0_root_sub_328_4_cf/U1_4  ( .A(n65606), .B(N11381), 
        .CI(\add_0_root_add_0_root_sub_328_4_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_328_4_cf/carry [5]), .S(N857) );
  ADD32 \add_0_root_add_0_root_sub_328_8_cf/U1_4  ( .A(N4178), .B(N11387), 
        .CI(\add_0_root_add_0_root_sub_328_8_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_328_8_cf/carry [5]), .S(N863) );
  ADD32 \add_0_root_add_0_root_sub_400_4_cf/U1_4  ( .A(n65608), .B(N11369), 
        .CI(\add_0_root_add_0_root_sub_400_4_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_400_4_cf/carry [5]), .S(N1145) );
  ADD32 \add_0_root_add_0_root_sub_400_8_cf/U1_4  ( .A(N6448), .B(N11375), 
        .CI(\add_0_root_add_0_root_sub_400_8_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_400_8_cf/carry [5]), .S(N1151) );
  ADD32 \add_0_root_add_0_root_sub_331_4_cf/U1_4  ( .A(n65608), .B(N11405), 
        .CI(\add_0_root_add_0_root_sub_331_4_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_331_4_cf/carry [5]), .S(N875) );
  ADD32 \add_0_root_add_0_root_sub_403_4_cf/U1_4  ( .A(n65606), .B(N11393), 
        .CI(\add_0_root_add_0_root_sub_403_4_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_403_4_cf/carry [5]), .S(N1163) );
  ADD32 \add_342_5/U1_4  ( .A(n65606), .B(n65597), .CI(\r38360/carry [4]), 
        .CO(\add_342_5/carry[5] ), .S(N941) );
  ADD32 \add_414_5/U1_4  ( .A(n65606), .B(n65597), .CI(\r38360/carry [4]), 
        .CO(\add_414_5/carry[5] ), .S(N1229) );
  ADD32 \add_345_3/U1_4  ( .A(n65607), .B(n65597), .CI(\r38360/carry [4]), 
        .CO(\add_345_3/carry[5] ), .S(N953) );
  ADD22 \sub_345_9_cf/U1_1_1  ( .A(n65758), .B(n65836), .CO(
        \sub_345_9_cf/carry [2]), .S(N956) );
  ADD22 \sub_345_9_cf/U1_1_2  ( .A(n65918), .B(\sub_345_9_cf/carry [2]), .CO(
        \sub_345_9_cf/carry [3]), .S(N957) );
  ADD22 \sub_345_9_cf/U1_1_3  ( .A(N11520), .B(\sub_345_9_cf/carry [3]), .CO(
        \sub_345_9_cf/carry [4]), .S(N958) );
  ADD22 \sub_345_9_cf/U1_1_4  ( .A(N11519), .B(\sub_345_9_cf/carry [4]), .CO(
        \sub_345_9_cf/carry [5]), .S(N959) );
  ADD32 \add_345_5/U1_4  ( .A(N4881), .B(n65599), .CI(\r32996/carry [4]), .CO(
        \add_345_5/carry[5] ), .S(N11519) );
  ADD32 \add_417_3/U1_4  ( .A(n65606), .B(n65598), .CI(\r38360/carry [4]), 
        .CO(\add_417_3/carry[5] ), .S(N1241) );
  ADD22 \sub_417_9_cf/U1_1_1  ( .A(n65758), .B(n65840), .CO(
        \sub_417_9_cf/carry [2]), .S(N1244) );
  ADD22 \sub_417_9_cf/U1_1_2  ( .A(n65918), .B(\sub_417_9_cf/carry [2]), .CO(
        \sub_417_9_cf/carry [3]), .S(N1245) );
  ADD22 \sub_417_9_cf/U1_1_3  ( .A(N11508), .B(\sub_417_9_cf/carry [3]), .CO(
        \sub_417_9_cf/carry [4]), .S(N1246) );
  ADD22 \sub_417_9_cf/U1_1_4  ( .A(N11507), .B(\sub_417_9_cf/carry [4]), .CO(
        \sub_417_9_cf/carry [5]), .S(N1247) );
  ADD32 \add_417_5/U1_4  ( .A(N7151), .B(n65597), .CI(\r32996/carry [4]), .CO(
        \add_417_5/carry[5] ), .S(N11507) );
  ADD32 \add_348/U1_4  ( .A(n65607), .B(n65598), .CI(\r38360/carry [4]), .CO(
        \add_348/carry[5] ), .S(N965) );
  ADD22 \sub_348_6_cf/U1_1_1  ( .A(n65758), .B(n65837), .CO(
        \sub_348_6_cf/carry [2]), .S(N968) );
  ADD22 \sub_348_6_cf/U1_1_2  ( .A(n65918), .B(\sub_348_6_cf/carry [2]), .CO(
        \sub_348_6_cf/carry [3]), .S(N969) );
  ADD22 \sub_348_6_cf/U1_1_3  ( .A(N11538), .B(\sub_348_6_cf/carry [3]), .CO(
        \sub_348_6_cf/carry [4]), .S(N970) );
  ADD22 \sub_348_6_cf/U1_1_4  ( .A(N11537), .B(\sub_348_6_cf/carry [4]), .CO(
        \sub_348_6_cf/carry [5]), .S(N971) );
  ADD32 \add_348_3/U1_4  ( .A(N5007), .B(n65597), .CI(\r32996/carry [4]), .CO(
        \add_348_3/carry[5] ), .S(N11537) );
  ADD32 \add_0_root_add_0_root_sub_348_9_cf/U1_4  ( .A(m[1]), .B(N11543), .CI(
        \add_0_root_add_0_root_sub_348_9_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_348_9_cf/carry [5]), .S(N977) );
  ADD32 \add_420/U1_4  ( .A(n65607), .B(n65597), .CI(\r38360/carry [4]), .CO(
        \add_420/carry[5] ), .S(N1253) );
  ADD22 \sub_420_6_cf/U1_1_1  ( .A(n65757), .B(n65838), .CO(
        \sub_420_6_cf/carry [2]), .S(N1256) );
  ADD22 \sub_420_6_cf/U1_1_2  ( .A(n65918), .B(\sub_420_6_cf/carry [2]), .CO(
        \sub_420_6_cf/carry [3]), .S(N1257) );
  ADD22 \sub_420_6_cf/U1_1_3  ( .A(N11526), .B(\sub_420_6_cf/carry [3]), .CO(
        \sub_420_6_cf/carry [4]), .S(N1258) );
  ADD22 \sub_420_6_cf/U1_1_4  ( .A(N11525), .B(\sub_420_6_cf/carry [4]), .CO(
        \sub_420_6_cf/carry [5]), .S(N1259) );
  ADD32 \add_420_3/U1_4  ( .A(N7277), .B(n65598), .CI(\r32996/carry [4]), .CO(
        \add_420_3/carry[5] ), .S(N11525) );
  ADD32 \add_0_root_add_0_root_sub_420_9_cf/U1_4  ( .A(m[1]), .B(N11531), .CI(
        \add_0_root_add_0_root_sub_420_9_cf/carry [4]), .CO(
        \add_0_root_add_0_root_sub_420_9_cf/carry [5]), .S(N1265) );
  ADD22 \add_1_root_add_126_3/U1_1_1  ( .A(G_play[1]), .B(n65532), .CO(
        \add_1_root_add_126_3/carry[2] ), .S(N1293) );
  ADD22 \add_1_root_add_126_3/U1_1_2  ( .A(G_play[2]), .B(
        \add_1_root_add_126_3/carry[2] ), .CO(N1295), .S(N1294) );
  ADD22 \r2195/U6  ( .A(N1836), .B(n65740), .CO(\r2195/n5 ), .S(N2049) );
  ADD32 \r2195/U5  ( .A(N1837), .B(N1836), .CI(\r2195/n5 ), .CO(\r2195/n4 ), 
        .S(N2050) );
  ADD32 \r2195/U4  ( .A(N1838), .B(N1837), .CI(\r2195/n4 ), .CO(\r2195/n3 ), 
        .S(N2051) );
  ADD22 \r2182/U6  ( .A(N1293), .B(n65742), .CO(\r2182/n5 ), .S(N1506) );
  ADD32 \r2182/U5  ( .A(N1294), .B(N1293), .CI(\r2182/n5 ), .CO(\r2182/n4 ), 
        .S(N1507) );
  ADD32 \r2182/U4  ( .A(N1295), .B(N1294), .CI(\r2182/n4 ), .CO(\r2182/n3 ), 
        .S(N1508) );
  ADD32 \r30599/U1_4  ( .A(N4593), .B(N11465), .CI(\r30599/carry [4]), .CO(
        \r30599/carry [5]), .S(N1205) );
  ADD32 \r30599/U1_5  ( .A(N4594), .B(N11464), .CI(\r30599/carry [5]), .S(
        N1206) );
  ADD22 \r31196/U1_1_2  ( .A(n65918), .B(\r31196/carry [2]), .CO(
        \r31196/carry [3]), .S(N1173) );
  ADD22 \r31196/U1_1_3  ( .A(N11412), .B(\r31196/carry [3]), .CO(
        \r31196/carry [4]), .S(N1174) );
  ADD22 \r31196/U1_1_4  ( .A(N11411), .B(\r31196/carry [4]), .CO(
        \r31196/carry [5]), .S(N1175) );
  ADD32 \r31195/U1_4  ( .A(N4329), .B(n65598), .CI(\r32996/carry [4]), .CO(
        \r31195/carry[5] ), .S(N11411) );
  ADD32 \r31798/U1_4  ( .A(N3204), .B(N3210), .CI(\r31798/carry [4]), .CO(
        \r31798/carry [5]), .S(N1019) );
  ADD32 \r31798/U1_5  ( .A(N3205), .B(N3211), .CI(\r31798/carry [5]), .S(N1020) );
  ADD32 \r32400/U1_4  ( .A(N3377), .B(N3383), .CI(\r32400/carry [4]), .CO(
        \r32400/carry [5]), .S(N1043) );
  ADD32 \r32400/U1_5  ( .A(N3378), .B(N3384), .CI(\r32400/carry [5]), .S(N1044) );
  ADD22 \r32997/U1_1_2  ( .A(n65918), .B(\r32997/carry [2]), .CO(
        \r32997/carry [3]), .S(N1185) );
  ADD22 \r32997/U1_1_3  ( .A(N11430), .B(\r32997/carry [3]), .CO(
        \r32997/carry [4]), .S(N1186) );
  ADD22 \r32997/U1_1_4  ( .A(N11429), .B(\r32997/carry [4]), .CO(
        \r32997/carry [5]), .S(N1187) );
  ADD32 \r32996/U1_4  ( .A(N4456), .B(n65597), .CI(\r32996/carry [4]), .CO(
        \r32996/carry [5]), .S(N11429) );
  ADD32 \r33599/U1_4  ( .A(N4730), .B(N11495), .CI(\r33599/carry [4]), .CO(
        \r33599/carry [5]), .S(N1223) );
  ADD32 \r33599/U1_5  ( .A(N4731), .B(N11494), .CI(\r33599/carry [5]), .S(
        N1224) );
  ADD32 \r34787/U1_4  ( .A(N4718), .B(N11489), .CI(\r34787/carry [4]), .CO(
        \r34787/carry [5]), .S(N1217) );
  ADD32 \r34787/U1_5  ( .A(N4719), .B(N11488), .CI(\r34787/carry [5]), .S(
        N1218) );
  ADD32 \r35376/U1_4  ( .A(N4444), .B(n65598), .CI(\r38360/carry [4]), .CO(
        \r35376/carry[5] ), .S(N1181) );
  ADD32 \r35376/U1_5  ( .A(N4445), .B(n[5]), .CI(\r35376/carry[5] ), .S(N1182)
         );
  ADD32 \r35965/U1_4  ( .A(N4190), .B(n[4]), .CI(\r38360/carry [4]), .CO(
        \r35965/carry[5] ), .S(N1157) );
  ADD32 \r35965/U1_5  ( .A(N4191), .B(n[5]), .CI(\r35965/carry[5] ), .S(N1158)
         );
  ADD32 \r36567/U1_4  ( .A(N3222), .B(N3228), .CI(\r36567/carry [4]), .CO(
        \r36567/carry [5]), .S(N1025) );
  ADD32 \r36567/U1_5  ( .A(N3223), .B(N3229), .CI(\r36567/carry [5]), .S(N1026) );
  ADD32 \r37169/U1_4  ( .A(N3049), .B(N3055), .CI(\r37169/carry [4]), .CO(
        \r37169/carry [5]), .S(N1001) );
  ADD32 \r37169/U1_5  ( .A(N3050), .B(N3056), .CI(\r37169/carry [5]), .S(N1002) );
  ADD32 \r37771/U1_4  ( .A(N3395), .B(N3401), .CI(\r37771/carry [4]), .CO(
        \r37771/carry [5]), .S(N1049) );
  ADD32 \r37771/U1_5  ( .A(N3396), .B(N3402), .CI(\r37771/carry [5]), .S(N1050) );
  ADD32 \r38360/U1_4  ( .A(N4317), .B(n65598), .CI(\r38360/carry [4]), .CO(
        \r38360/carry [5]), .S(N1169) );
  ADD32 \r38360/U1_5  ( .A(N4318), .B(n65600), .CI(\r38360/carry [5]), .S(
        N1170) );
  ADD32 \r38962/U1_4  ( .A(N4581), .B(N11459), .CI(\r38962/carry [4]), .CO(
        \r38962/carry [5]), .S(N1199) );
  ADD32 \r38962/U1_5  ( .A(N4582), .B(N11458), .CI(\r38962/carry [5]), .S(
        N1200) );
  ADD32 \r39564/U1_4  ( .A(N4857), .B(N11513), .CI(\r39564/carry [4]), .CO(
        \r39564/carry [5]), .S(N1235) );
  ADD32 \r39564/U1_5  ( .A(N4858), .B(N11512), .CI(\r39564/carry [5]), .S(
        N1236) );
  ADD32 \r40166/U1_4  ( .A(N4468), .B(N11435), .CI(\r40166/carry [4]), .CO(
        \r40166/carry [5]), .S(N1193) );
  ADD32 \r40166/U1_5  ( .A(N4469), .B(N11434), .CI(\r40166/carry [5]), .S(
        N1194) );
  ADD32 \r40768/U1_4  ( .A(N3359), .B(N3365), .CI(\r40768/carry [4]), .CO(
        \r40768/carry [5]), .S(N1037) );
  ADD32 \r40768/U1_5  ( .A(N3360), .B(N3366), .CI(\r40768/carry [5]), .S(N1038) );
  ADD32 \r41370/U1_4  ( .A(N4605), .B(N11471), .CI(\r41370/carry [4]), .CO(
        \r41370/carry [5]), .S(N1211) );
  ADD32 \r41370/U1_5  ( .A(N4606), .B(N11470), .CI(\r41370/carry [5]), .S(
        N1212) );
  IMUX40 U7553 ( .A(\Col_Fill[0][29] ), .B(\Col_Fill[1][29] ), .C(
        \Col_Fill[2][29] ), .D(\Col_Fill[3][29] ), .S0(n65512), .S1(N689), .Q(
        n3973) );
  IMUX40 U7552 ( .A(\Col_Fill[4][29] ), .B(\Col_Fill[5][29] ), .C(
        \Col_Fill[6][29] ), .D(\Col_Fill[7][29] ), .S0(n65522), .S1(n65939), 
        .Q(n3974) );
  IMUX21 U7491 ( .A(n3973), .B(n3974), .S(n65937), .Q(N1984) );
  IMUX40 U7361 ( .A(\Col_Fill[0][29] ), .B(\Col_Fill[1][29] ), .C(
        \Col_Fill[2][29] ), .D(\Col_Fill[3][29] ), .S0(n65533), .S1(N683), .Q(
        n3845) );
  IMUX40 U7360 ( .A(\Col_Fill[4][29] ), .B(\Col_Fill[5][29] ), .C(
        \Col_Fill[6][29] ), .D(\Col_Fill[7][29] ), .S0(n65532), .S1(n65949), 
        .Q(n3846) );
  IMUX21 U7299 ( .A(n3845), .B(n3846), .S(n65947), .Q(N1441) );
  IMUX40 U7551 ( .A(\Col_Fill[0][28] ), .B(\Col_Fill[1][28] ), .C(
        \Col_Fill[2][28] ), .D(\Col_Fill[3][28] ), .S0(n65511), .S1(n65938), 
        .Q(n3971) );
  IMUX40 U7550 ( .A(\Col_Fill[4][28] ), .B(\Col_Fill[5][28] ), .C(
        \Col_Fill[6][28] ), .D(\Col_Fill[7][28] ), .S0(n65522), .S1(n65941), 
        .Q(n3972) );
  IMUX21 U7490 ( .A(n3971), .B(n3972), .S(n65937), .Q(N1985) );
  IMUX40 U7359 ( .A(\Col_Fill[0][28] ), .B(\Col_Fill[1][28] ), .C(
        \Col_Fill[2][28] ), .D(\Col_Fill[3][28] ), .S0(n65533), .S1(n65948), 
        .Q(n3843) );
  IMUX40 U7358 ( .A(\Col_Fill[4][28] ), .B(\Col_Fill[5][28] ), .C(
        \Col_Fill[6][28] ), .D(\Col_Fill[7][28] ), .S0(n65532), .S1(n65951), 
        .Q(n3844) );
  IMUX21 U7298 ( .A(n3843), .B(n3844), .S(n65947), .Q(N1442) );
  IMUX40 U7549 ( .A(\Col_Fill[0][27] ), .B(\Col_Fill[1][27] ), .C(
        \Col_Fill[2][27] ), .D(\Col_Fill[3][27] ), .S0(n65520), .S1(n65939), 
        .Q(n3969) );
  IMUX40 U7548 ( .A(\Col_Fill[4][27] ), .B(\Col_Fill[5][27] ), .C(
        \Col_Fill[6][27] ), .D(\Col_Fill[7][27] ), .S0(n65520), .S1(n65940), 
        .Q(n3970) );
  IMUX21 U7489 ( .A(n3969), .B(n3970), .S(N690), .Q(N1986) );
  IMUX40 U7357 ( .A(\Col_Fill[0][27] ), .B(\Col_Fill[1][27] ), .C(
        \Col_Fill[2][27] ), .D(\Col_Fill[3][27] ), .S0(n65420), .S1(n65949), 
        .Q(n3841) );
  IMUX40 U7356 ( .A(\Col_Fill[4][27] ), .B(\Col_Fill[5][27] ), .C(
        \Col_Fill[6][27] ), .D(\Col_Fill[7][27] ), .S0(n65530), .S1(n65950), 
        .Q(n3842) );
  IMUX21 U7297 ( .A(n3841), .B(n3842), .S(N684), .Q(N1443) );
  IMUX40 U7547 ( .A(\Col_Fill[0][26] ), .B(\Col_Fill[1][26] ), .C(
        \Col_Fill[2][26] ), .D(\Col_Fill[3][26] ), .S0(n65521), .S1(n65941), 
        .Q(n3967) );
  IMUX40 U7546 ( .A(\Col_Fill[4][26] ), .B(\Col_Fill[5][26] ), .C(
        \Col_Fill[6][26] ), .D(\Col_Fill[7][26] ), .S0(n65520), .S1(N689), .Q(
        n3968) );
  IMUX21 U7488 ( .A(n3967), .B(n3968), .S(n65937), .Q(N1987) );
  IMUX40 U7355 ( .A(\Col_Fill[0][26] ), .B(\Col_Fill[1][26] ), .C(
        \Col_Fill[2][26] ), .D(\Col_Fill[3][26] ), .S0(n65527), .S1(n65951), 
        .Q(n3839) );
  IMUX40 U7354 ( .A(\Col_Fill[4][26] ), .B(\Col_Fill[5][26] ), .C(
        \Col_Fill[6][26] ), .D(\Col_Fill[7][26] ), .S0(n65524), .S1(N683), .Q(
        n3840) );
  IMUX21 U7296 ( .A(n3839), .B(n3840), .S(n65947), .Q(N1444) );
  IMUX40 U7545 ( .A(\Col_Fill[0][25] ), .B(\Col_Fill[1][25] ), .C(
        \Col_Fill[2][25] ), .D(\Col_Fill[3][25] ), .S0(n65514), .S1(n65942), 
        .Q(n3965) );
  IMUX40 U7544 ( .A(\Col_Fill[4][25] ), .B(\Col_Fill[5][25] ), .C(
        \Col_Fill[6][25] ), .D(\Col_Fill[7][25] ), .S0(n65521), .S1(n65945), 
        .Q(n3966) );
  IMUX21 U7487 ( .A(n3965), .B(n3966), .S(N690), .Q(N1988) );
  IMUX40 U7353 ( .A(\Col_Fill[0][25] ), .B(\Col_Fill[1][25] ), .C(
        \Col_Fill[2][25] ), .D(\Col_Fill[3][25] ), .S0(n65528), .S1(n65952), 
        .Q(n3837) );
  IMUX40 U7352 ( .A(\Col_Fill[4][25] ), .B(\Col_Fill[5][25] ), .C(
        \Col_Fill[6][25] ), .D(\Col_Fill[7][25] ), .S0(n65525), .S1(n65955), 
        .Q(n3838) );
  IMUX21 U7295 ( .A(n3837), .B(n3838), .S(N684), .Q(N1445) );
  IMUX40 U7543 ( .A(\Col_Fill[0][24] ), .B(\Col_Fill[1][24] ), .C(
        \Col_Fill[2][24] ), .D(\Col_Fill[3][24] ), .S0(n65520), .S1(n65944), 
        .Q(n3963) );
  IMUX40 U7542 ( .A(\Col_Fill[4][24] ), .B(\Col_Fill[5][24] ), .C(
        \Col_Fill[6][24] ), .D(\Col_Fill[7][24] ), .S0(n65514), .S1(n65941), 
        .Q(n3964) );
  IMUX21 U7486 ( .A(n3963), .B(n3964), .S(n65937), .Q(N1989) );
  IMUX40 U7351 ( .A(\Col_Fill[0][24] ), .B(\Col_Fill[1][24] ), .C(
        \Col_Fill[2][24] ), .D(\Col_Fill[3][24] ), .S0(n65531), .S1(n65951), 
        .Q(n3835) );
  IMUX40 U7350 ( .A(\Col_Fill[4][24] ), .B(\Col_Fill[5][24] ), .C(
        \Col_Fill[6][24] ), .D(\Col_Fill[7][24] ), .S0(n65533), .S1(n65954), 
        .Q(n3836) );
  IMUX21 U7294 ( .A(n3835), .B(n3836), .S(n65947), .Q(N1446) );
  IMUX40 U7541 ( .A(\Col_Fill[0][23] ), .B(\Col_Fill[1][23] ), .C(
        \Col_Fill[2][23] ), .D(\Col_Fill[3][23] ), .S0(n65521), .S1(n65943), 
        .Q(n3961) );
  IMUX40 U7540 ( .A(\Col_Fill[4][23] ), .B(\Col_Fill[5][23] ), .C(
        \Col_Fill[6][23] ), .D(\Col_Fill[7][23] ), .S0(n65520), .S1(n65939), 
        .Q(n3962) );
  IMUX21 U7485 ( .A(n3961), .B(n3962), .S(N690), .Q(N1990) );
  IMUX40 U7349 ( .A(\Col_Fill[0][23] ), .B(\Col_Fill[1][23] ), .C(
        \Col_Fill[2][23] ), .D(\Col_Fill[3][23] ), .S0(n65453), .S1(n65953), 
        .Q(n3833) );
  IMUX40 U7348 ( .A(\Col_Fill[4][23] ), .B(\Col_Fill[5][23] ), .C(
        \Col_Fill[6][23] ), .D(\Col_Fill[7][23] ), .S0(n65453), .S1(n65949), 
        .Q(n3834) );
  IMUX21 U7293 ( .A(n3833), .B(n3834), .S(N684), .Q(N1447) );
  IMUX40 U7539 ( .A(\Col_Fill[0][22] ), .B(\Col_Fill[1][22] ), .C(
        \Col_Fill[2][22] ), .D(\Col_Fill[3][22] ), .S0(n65515), .S1(n65938), 
        .Q(n3959) );
  IMUX40 U7538 ( .A(\Col_Fill[4][22] ), .B(\Col_Fill[5][22] ), .C(
        \Col_Fill[6][22] ), .D(\Col_Fill[7][22] ), .S0(n65521), .S1(n65941), 
        .Q(n3960) );
  IMUX21 U7484 ( .A(n3959), .B(n3960), .S(n65937), .Q(N1991) );
  IMUX40 U7347 ( .A(\Col_Fill[0][22] ), .B(\Col_Fill[1][22] ), .C(
        \Col_Fill[2][22] ), .D(\Col_Fill[3][22] ), .S0(n65526), .S1(n65948), 
        .Q(n3831) );
  IMUX40 U7346 ( .A(\Col_Fill[4][22] ), .B(\Col_Fill[5][22] ), .C(
        \Col_Fill[6][22] ), .D(\Col_Fill[7][22] ), .S0(n65529), .S1(n65951), 
        .Q(n3832) );
  IMUX21 U7292 ( .A(n3831), .B(n3832), .S(n65947), .Q(N1448) );
  IMUX40 U7537 ( .A(\Col_Fill[0][21] ), .B(\Col_Fill[1][21] ), .C(
        \Col_Fill[2][21] ), .D(\Col_Fill[3][21] ), .S0(n65514), .S1(n65939), 
        .Q(n3957) );
  IMUX40 U7536 ( .A(\Col_Fill[4][21] ), .B(\Col_Fill[5][21] ), .C(
        \Col_Fill[6][21] ), .D(\Col_Fill[7][21] ), .S0(n65518), .S1(n65940), 
        .Q(n3958) );
  IMUX21 U7483 ( .A(n3957), .B(n3958), .S(N690), .Q(N1992) );
  IMUX40 U7345 ( .A(\Col_Fill[0][21] ), .B(\Col_Fill[1][21] ), .C(
        \Col_Fill[2][21] ), .D(\Col_Fill[3][21] ), .S0(n65526), .S1(n65949), 
        .Q(n3829) );
  IMUX40 U7344 ( .A(\Col_Fill[4][21] ), .B(\Col_Fill[5][21] ), .C(
        \Col_Fill[6][21] ), .D(\Col_Fill[7][21] ), .S0(n65420), .S1(n65950), 
        .Q(n3830) );
  IMUX21 U7291 ( .A(n3829), .B(n3830), .S(N684), .Q(N1449) );
  IMUX40 U7535 ( .A(\Col_Fill[0][20] ), .B(\Col_Fill[1][20] ), .C(
        \Col_Fill[2][20] ), .D(\Col_Fill[3][20] ), .S0(n65519), .S1(n65938), 
        .Q(n3955) );
  IMUX40 U7534 ( .A(\Col_Fill[4][20] ), .B(\Col_Fill[5][20] ), .C(
        \Col_Fill[6][20] ), .D(\Col_Fill[7][20] ), .S0(n65519), .S1(n65945), 
        .Q(n3956) );
  IMUX21 U7482 ( .A(n3955), .B(n3956), .S(n65937), .Q(N1993) );
  IMUX40 U7343 ( .A(\Col_Fill[0][20] ), .B(\Col_Fill[1][20] ), .C(
        \Col_Fill[2][20] ), .D(\Col_Fill[3][20] ), .S0(n65524), .S1(n65948), 
        .Q(n3827) );
  IMUX40 U7342 ( .A(\Col_Fill[4][20] ), .B(\Col_Fill[5][20] ), .C(
        \Col_Fill[6][20] ), .D(\Col_Fill[7][20] ), .S0(n65420), .S1(n65955), 
        .Q(n3828) );
  IMUX21 U7290 ( .A(n3827), .B(n3828), .S(n65947), .Q(N1450) );
  IMUX40 U7533 ( .A(\Col_Fill[0][19] ), .B(\Col_Fill[1][19] ), .C(
        \Col_Fill[2][19] ), .D(\Col_Fill[3][19] ), .S0(n65518), .S1(n65942), 
        .Q(n3953) );
  IMUX40 U7532 ( .A(\Col_Fill[4][19] ), .B(\Col_Fill[5][19] ), .C(
        \Col_Fill[6][19] ), .D(\Col_Fill[7][19] ), .S0(n65519), .S1(n65942), 
        .Q(n3954) );
  IMUX21 U7481 ( .A(n3953), .B(n3954), .S(N690), .Q(N1994) );
  IMUX40 U7341 ( .A(\Col_Fill[0][19] ), .B(\Col_Fill[1][19] ), .C(
        \Col_Fill[2][19] ), .D(\Col_Fill[3][19] ), .S0(n65420), .S1(n65952), 
        .Q(n3825) );
  IMUX40 U7340 ( .A(\Col_Fill[4][19] ), .B(\Col_Fill[5][19] ), .C(
        \Col_Fill[6][19] ), .D(\Col_Fill[7][19] ), .S0(n65453), .S1(n65952), 
        .Q(n3826) );
  IMUX21 U7289 ( .A(n3825), .B(n3826), .S(N684), .Q(N1451) );
  IMUX40 U7531 ( .A(\Col_Fill[0][18] ), .B(\Col_Fill[1][18] ), .C(
        \Col_Fill[2][18] ), .D(\Col_Fill[3][18] ), .S0(n65419), .S1(n65942), 
        .Q(n3951) );
  IMUX40 U7530 ( .A(\Col_Fill[4][18] ), .B(\Col_Fill[5][18] ), .C(
        \Col_Fill[6][18] ), .D(\Col_Fill[7][18] ), .S0(n65518), .S1(n65942), 
        .Q(n3952) );
  IMUX21 U7480 ( .A(n3951), .B(n3952), .S(n65937), .Q(N1995) );
  IMUX40 U7339 ( .A(\Col_Fill[0][18] ), .B(\Col_Fill[1][18] ), .C(
        \Col_Fill[2][18] ), .D(\Col_Fill[3][18] ), .S0(n65453), .S1(n65952), 
        .Q(n3823) );
  IMUX40 U7338 ( .A(\Col_Fill[4][18] ), .B(\Col_Fill[5][18] ), .C(
        \Col_Fill[6][18] ), .D(\Col_Fill[7][18] ), .S0(n65453), .S1(n65952), 
        .Q(n3824) );
  IMUX21 U7288 ( .A(n3823), .B(n3824), .S(n65947), .Q(N1452) );
  IMUX40 U7529 ( .A(\Col_Fill[0][17] ), .B(\Col_Fill[1][17] ), .C(
        \Col_Fill[2][17] ), .D(\Col_Fill[3][17] ), .S0(n65519), .S1(n65942), 
        .Q(n3949) );
  IMUX40 U7528 ( .A(\Col_Fill[4][17] ), .B(\Col_Fill[5][17] ), .C(
        \Col_Fill[6][17] ), .D(\Col_Fill[7][17] ), .S0(n65511), .S1(n65942), 
        .Q(n3950) );
  IMUX21 U7479 ( .A(n3949), .B(n3950), .S(N690), .Q(N1996) );
  IMUX40 U7337 ( .A(\Col_Fill[0][17] ), .B(\Col_Fill[1][17] ), .C(
        \Col_Fill[2][17] ), .D(\Col_Fill[3][17] ), .S0(n65530), .S1(n65952), 
        .Q(n3821) );
  IMUX40 U7336 ( .A(\Col_Fill[4][17] ), .B(\Col_Fill[5][17] ), .C(
        \Col_Fill[6][17] ), .D(\Col_Fill[7][17] ), .S0(n65528), .S1(n65952), 
        .Q(n3822) );
  IMUX21 U7287 ( .A(n3821), .B(n3822), .S(N684), .Q(N1453) );
  IMUX40 U7527 ( .A(\Col_Fill[0][16] ), .B(\Col_Fill[1][16] ), .C(
        \Col_Fill[2][16] ), .D(\Col_Fill[3][16] ), .S0(n65518), .S1(n65942), 
        .Q(n3947) );
  IMUX40 U7526 ( .A(\Col_Fill[4][16] ), .B(\Col_Fill[5][16] ), .C(
        \Col_Fill[6][16] ), .D(\Col_Fill[7][16] ), .S0(n65519), .S1(n65942), 
        .Q(n3948) );
  IMUX21 U7478 ( .A(n3947), .B(n3948), .S(N690), .Q(N1997) );
  IMUX40 U7335 ( .A(\Col_Fill[0][16] ), .B(\Col_Fill[1][16] ), .C(
        \Col_Fill[2][16] ), .D(\Col_Fill[3][16] ), .S0(n65453), .S1(n65952), 
        .Q(n3819) );
  IMUX40 U7334 ( .A(\Col_Fill[4][16] ), .B(\Col_Fill[5][16] ), .C(
        \Col_Fill[6][16] ), .D(\Col_Fill[7][16] ), .S0(n65420), .S1(n65952), 
        .Q(n3820) );
  IMUX21 U7286 ( .A(n3819), .B(n3820), .S(N684), .Q(N1454) );
  IMUX40 U7525 ( .A(\Col_Fill[0][15] ), .B(\Col_Fill[1][15] ), .C(
        \Col_Fill[2][15] ), .D(\Col_Fill[3][15] ), .S0(n65511), .S1(n65942), 
        .Q(n3945) );
  IMUX40 U7524 ( .A(\Col_Fill[4][15] ), .B(\Col_Fill[5][15] ), .C(
        \Col_Fill[6][15] ), .D(\Col_Fill[7][15] ), .S0(n65521), .S1(n65942), 
        .Q(n3946) );
  IMUX21 U7477 ( .A(n3945), .B(n3946), .S(n65937), .Q(N1998) );
  IMUX40 U7333 ( .A(\Col_Fill[0][15] ), .B(\Col_Fill[1][15] ), .C(
        \Col_Fill[2][15] ), .D(\Col_Fill[3][15] ), .S0(n65420), .S1(n65952), 
        .Q(n3817) );
  IMUX40 U7332 ( .A(\Col_Fill[4][15] ), .B(\Col_Fill[5][15] ), .C(
        \Col_Fill[6][15] ), .D(\Col_Fill[7][15] ), .S0(n65532), .S1(n65952), 
        .Q(n3818) );
  IMUX21 U7285 ( .A(n3817), .B(n3818), .S(n65946), .Q(N1455) );
  IMUX40 U7523 ( .A(\Col_Fill[0][14] ), .B(\Col_Fill[1][14] ), .C(
        \Col_Fill[2][14] ), .D(\Col_Fill[3][14] ), .S0(n65516), .S1(n65942), 
        .Q(n3943) );
  IMUX40 U7522 ( .A(\Col_Fill[4][14] ), .B(\Col_Fill[5][14] ), .C(
        \Col_Fill[6][14] ), .D(\Col_Fill[7][14] ), .S0(n65522), .S1(n65942), 
        .Q(n3944) );
  IMUX21 U7476 ( .A(n3943), .B(n3944), .S(n65936), .Q(N1999) );
  IMUX40 U7331 ( .A(\Col_Fill[0][14] ), .B(\Col_Fill[1][14] ), .C(
        \Col_Fill[2][14] ), .D(\Col_Fill[3][14] ), .S0(n65523), .S1(n65952), 
        .Q(n3815) );
  IMUX40 U7330 ( .A(\Col_Fill[4][14] ), .B(\Col_Fill[5][14] ), .C(
        \Col_Fill[6][14] ), .D(\Col_Fill[7][14] ), .S0(n65524), .S1(n65952), 
        .Q(n3816) );
  IMUX21 U7284 ( .A(n3815), .B(n3816), .S(n65947), .Q(N1456) );
  IMUX40 U7521 ( .A(\Col_Fill[0][13] ), .B(\Col_Fill[1][13] ), .C(
        \Col_Fill[2][13] ), .D(\Col_Fill[3][13] ), .S0(n65510), .S1(n65940), 
        .Q(n3941) );
  IMUX40 U7520 ( .A(\Col_Fill[4][13] ), .B(\Col_Fill[5][13] ), .C(
        \Col_Fill[6][13] ), .D(\Col_Fill[7][13] ), .S0(n65522), .S1(n65941), 
        .Q(n3942) );
  IMUX21 U7475 ( .A(n3941), .B(n3942), .S(N690), .Q(N2000) );
  IMUX40 U7329 ( .A(\Col_Fill[0][13] ), .B(\Col_Fill[1][13] ), .C(
        \Col_Fill[2][13] ), .D(\Col_Fill[3][13] ), .S0(n65531), .S1(n65950), 
        .Q(n3813) );
  IMUX40 U7328 ( .A(\Col_Fill[4][13] ), .B(\Col_Fill[5][13] ), .C(
        \Col_Fill[6][13] ), .D(\Col_Fill[7][13] ), .S0(n65526), .S1(n65951), 
        .Q(n3814) );
  IMUX21 U7283 ( .A(n3813), .B(n3814), .S(N684), .Q(N1457) );
  IMUX40 U7519 ( .A(\Col_Fill[0][12] ), .B(\Col_Fill[1][12] ), .C(
        \Col_Fill[2][12] ), .D(\Col_Fill[3][12] ), .S0(n65515), .S1(n65939), 
        .Q(n3939) );
  IMUX40 U7518 ( .A(\Col_Fill[4][12] ), .B(\Col_Fill[5][12] ), .C(
        \Col_Fill[6][12] ), .D(\Col_Fill[7][12] ), .S0(n65520), .S1(n65938), 
        .Q(n3940) );
  IMUX21 U7474 ( .A(n3939), .B(n3940), .S(n65937), .Q(N2001) );
  IMUX40 U7327 ( .A(\Col_Fill[0][12] ), .B(\Col_Fill[1][12] ), .C(
        \Col_Fill[2][12] ), .D(\Col_Fill[3][12] ), .S0(n65533), .S1(n65949), 
        .Q(n3811) );
  IMUX40 U7326 ( .A(\Col_Fill[4][12] ), .B(\Col_Fill[5][12] ), .C(
        \Col_Fill[6][12] ), .D(\Col_Fill[7][12] ), .S0(n65420), .S1(n65948), 
        .Q(n3812) );
  IMUX21 U7282 ( .A(n3811), .B(n3812), .S(n65947), .Q(N1458) );
  IMUX40 U7517 ( .A(\Col_Fill[0][11] ), .B(\Col_Fill[1][11] ), .C(
        \Col_Fill[2][11] ), .D(\Col_Fill[3][11] ), .S0(n65511), .S1(n65941), 
        .Q(n3937) );
  IMUX40 U7516 ( .A(\Col_Fill[4][11] ), .B(\Col_Fill[5][11] ), .C(
        \Col_Fill[6][11] ), .D(\Col_Fill[7][11] ), .S0(n65517), .S1(n65945), 
        .Q(n3938) );
  IMUX21 U7473 ( .A(n3937), .B(n3938), .S(N690), .Q(N2002) );
  IMUX40 U7325 ( .A(\Col_Fill[0][11] ), .B(\Col_Fill[1][11] ), .C(
        \Col_Fill[2][11] ), .D(\Col_Fill[3][11] ), .S0(n65527), .S1(n65951), 
        .Q(n3809) );
  IMUX40 U7324 ( .A(\Col_Fill[4][11] ), .B(\Col_Fill[5][11] ), .C(
        \Col_Fill[6][11] ), .D(\Col_Fill[7][11] ), .S0(n65453), .S1(n65955), 
        .Q(n3810) );
  IMUX21 U7281 ( .A(n3809), .B(n3810), .S(n65946), .Q(N1459) );
  IMUX40 U7515 ( .A(\Col_Fill[0][10] ), .B(\Col_Fill[1][10] ), .C(
        \Col_Fill[2][10] ), .D(\Col_Fill[3][10] ), .S0(n65516), .S1(n65938), 
        .Q(n3935) );
  IMUX40 U7514 ( .A(\Col_Fill[4][10] ), .B(\Col_Fill[5][10] ), .C(
        \Col_Fill[6][10] ), .D(\Col_Fill[7][10] ), .S0(n65521), .S1(n65940), 
        .Q(n3936) );
  IMUX21 U7472 ( .A(n3935), .B(n3936), .S(n65936), .Q(N2003) );
  IMUX40 U7323 ( .A(\Col_Fill[0][10] ), .B(\Col_Fill[1][10] ), .C(
        \Col_Fill[2][10] ), .D(\Col_Fill[3][10] ), .S0(n65524), .S1(n65948), 
        .Q(n3807) );
  IMUX40 U7322 ( .A(\Col_Fill[4][10] ), .B(\Col_Fill[5][10] ), .C(
        \Col_Fill[6][10] ), .D(\Col_Fill[7][10] ), .S0(n65525), .S1(n65950), 
        .Q(n3808) );
  IMUX21 U7280 ( .A(n3807), .B(n3808), .S(N684), .Q(N1460) );
  IMUX40 U7513 ( .A(\Col_Fill[0][9] ), .B(\Col_Fill[1][9] ), .C(
        \Col_Fill[2][9] ), .D(\Col_Fill[3][9] ), .S0(n65419), .S1(n65945), .Q(
        n3933) );
  IMUX40 U7512 ( .A(\Col_Fill[4][9] ), .B(\Col_Fill[5][9] ), .C(
        \Col_Fill[6][9] ), .D(\Col_Fill[7][9] ), .S0(n65512), .S1(n65939), .Q(
        n3934) );
  IMUX21 U7471 ( .A(n3933), .B(n3934), .S(N690), .Q(N2004) );
  IMUX40 U7321 ( .A(\Col_Fill[0][9] ), .B(\Col_Fill[1][9] ), .C(
        \Col_Fill[2][9] ), .D(\Col_Fill[3][9] ), .S0(n65528), .S1(n65955), .Q(
        n3805) );
  IMUX40 U7320 ( .A(\Col_Fill[4][9] ), .B(\Col_Fill[5][9] ), .C(
        \Col_Fill[6][9] ), .D(\Col_Fill[7][9] ), .S0(n65529), .S1(n65949), .Q(
        n3806) );
  IMUX21 U7279 ( .A(n3805), .B(n3806), .S(N684), .Q(N1461) );
  IMUX40 U7511 ( .A(\Col_Fill[0][8] ), .B(\Col_Fill[1][8] ), .C(
        \Col_Fill[2][8] ), .D(\Col_Fill[3][8] ), .S0(n65519), .S1(n65939), .Q(
        n3931) );
  IMUX40 U7510 ( .A(\Col_Fill[4][8] ), .B(\Col_Fill[5][8] ), .C(
        \Col_Fill[6][8] ), .D(\Col_Fill[7][8] ), .S0(n65419), .S1(n65941), .Q(
        n3932) );
  IMUX21 U7470 ( .A(n3931), .B(n3932), .S(n65937), .Q(N2005) );
  IMUX40 U7319 ( .A(\Col_Fill[0][8] ), .B(\Col_Fill[1][8] ), .C(
        \Col_Fill[2][8] ), .D(\Col_Fill[3][8] ), .S0(n65530), .S1(n65949), .Q(
        n3803) );
  IMUX40 U7318 ( .A(\Col_Fill[4][8] ), .B(\Col_Fill[5][8] ), .C(
        \Col_Fill[6][8] ), .D(\Col_Fill[7][8] ), .S0(n65528), .S1(n65951), .Q(
        n3804) );
  IMUX21 U7278 ( .A(n3803), .B(n3804), .S(n65947), .Q(N1462) );
  IMUX40 U7509 ( .A(\Col_Fill[0][7] ), .B(\Col_Fill[1][7] ), .C(
        \Col_Fill[2][7] ), .D(\Col_Fill[3][7] ), .S0(n65419), .S1(n65939), .Q(
        n3929) );
  IMUX40 U7508 ( .A(\Col_Fill[4][7] ), .B(\Col_Fill[5][7] ), .C(
        \Col_Fill[6][7] ), .D(\Col_Fill[7][7] ), .S0(n65512), .S1(n65938), .Q(
        n3930) );
  IMUX21 U7469 ( .A(n3929), .B(n3930), .S(N690), .Q(N2006) );
  IMUX40 U7317 ( .A(\Col_Fill[0][7] ), .B(\Col_Fill[1][7] ), .C(
        \Col_Fill[2][7] ), .D(\Col_Fill[3][7] ), .S0(n65529), .S1(n65949), .Q(
        n3801) );
  IMUX40 U7316 ( .A(\Col_Fill[4][7] ), .B(\Col_Fill[5][7] ), .C(
        \Col_Fill[6][7] ), .D(\Col_Fill[7][7] ), .S0(n65530), .S1(n65948), .Q(
        n3802) );
  IMUX21 U7277 ( .A(n3801), .B(n3802), .S(N684), .Q(N1463) );
  IMUX40 U7507 ( .A(\Col_Fill[0][6] ), .B(\Col_Fill[1][6] ), .C(
        \Col_Fill[2][6] ), .D(\Col_Fill[3][6] ), .S0(n65419), .S1(n65945), .Q(
        n3927) );
  IMUX40 U7506 ( .A(\Col_Fill[4][6] ), .B(\Col_Fill[5][6] ), .C(
        \Col_Fill[6][6] ), .D(\Col_Fill[7][6] ), .S0(n65518), .S1(n65940), .Q(
        n3928) );
  IMUX21 U7468 ( .A(n3927), .B(n3928), .S(n65937), .Q(N2007) );
  IMUX40 U7315 ( .A(\Col_Fill[0][6] ), .B(\Col_Fill[1][6] ), .C(
        \Col_Fill[2][6] ), .D(\Col_Fill[3][6] ), .S0(n65528), .S1(n65955), .Q(
        n3799) );
  IMUX40 U7314 ( .A(\Col_Fill[4][6] ), .B(\Col_Fill[5][6] ), .C(
        \Col_Fill[6][6] ), .D(\Col_Fill[7][6] ), .S0(n65529), .S1(n65950), .Q(
        n3800) );
  IMUX21 U7276 ( .A(n3799), .B(n3800), .S(n65947), .Q(N1464) );
  IMUX40 U7505 ( .A(\Col_Fill[0][5] ), .B(\Col_Fill[1][5] ), .C(
        \Col_Fill[2][5] ), .D(\Col_Fill[3][5] ), .S0(n65520), .S1(n65940), .Q(
        n3925) );
  IMUX40 U7504 ( .A(\Col_Fill[4][5] ), .B(\Col_Fill[5][5] ), .C(
        \Col_Fill[6][5] ), .D(\Col_Fill[7][5] ), .S0(n65518), .S1(n65943), .Q(
        n3926) );
  IMUX21 U7467 ( .A(n3925), .B(n3926), .S(N690), .Q(N2008) );
  IMUX40 U7313 ( .A(\Col_Fill[0][5] ), .B(\Col_Fill[1][5] ), .C(
        \Col_Fill[2][5] ), .D(\Col_Fill[3][5] ), .S0(n65530), .S1(n65954), .Q(
        n3797) );
  IMUX40 U7312 ( .A(\Col_Fill[4][5] ), .B(\Col_Fill[5][5] ), .C(
        \Col_Fill[6][5] ), .D(\Col_Fill[7][5] ), .S0(n65528), .S1(n65953), .Q(
        n3798) );
  IMUX21 U7275 ( .A(n3797), .B(n3798), .S(N684), .Q(N1465) );
  IMUX40 U7503 ( .A(\Col_Fill[0][4] ), .B(\Col_Fill[1][4] ), .C(
        \Col_Fill[2][4] ), .D(\Col_Fill[3][4] ), .S0(n65519), .S1(n65942), .Q(
        n3923) );
  IMUX40 U7502 ( .A(\Col_Fill[4][4] ), .B(\Col_Fill[5][4] ), .C(
        \Col_Fill[6][4] ), .D(\Col_Fill[7][4] ), .S0(n65510), .S1(n65944), .Q(
        n3924) );
  IMUX21 U7466 ( .A(n3923), .B(n3924), .S(n65937), .Q(N2009) );
  IMUX40 U7311 ( .A(\Col_Fill[0][4] ), .B(\Col_Fill[1][4] ), .C(
        \Col_Fill[2][4] ), .D(\Col_Fill[3][4] ), .S0(n65529), .S1(n65952), .Q(
        n3795) );
  IMUX40 U7310 ( .A(\Col_Fill[4][4] ), .B(\Col_Fill[5][4] ), .C(
        \Col_Fill[6][4] ), .D(\Col_Fill[7][4] ), .S0(n65530), .S1(n65950), .Q(
        n3796) );
  IMUX21 U7274 ( .A(n3795), .B(n3796), .S(n65947), .Q(N1466) );
  IMUX40 U7501 ( .A(\Col_Fill[0][3] ), .B(\Col_Fill[1][3] ), .C(
        \Col_Fill[2][3] ), .D(\Col_Fill[3][3] ), .S0(n65516), .S1(n65938), .Q(
        n3921) );
  IMUX40 U7500 ( .A(\Col_Fill[4][3] ), .B(\Col_Fill[5][3] ), .C(
        \Col_Fill[6][3] ), .D(\Col_Fill[7][3] ), .S0(n65419), .S1(n65941), .Q(
        n3922) );
  IMUX21 U7465 ( .A(n3921), .B(n3922), .S(n65936), .Q(N2010) );
  IMUX40 U7309 ( .A(\Col_Fill[0][3] ), .B(\Col_Fill[1][3] ), .C(
        \Col_Fill[2][3] ), .D(\Col_Fill[3][3] ), .S0(n65453), .S1(n65948), .Q(
        n3793) );
  IMUX40 U7308 ( .A(\Col_Fill[4][3] ), .B(\Col_Fill[5][3] ), .C(
        \Col_Fill[6][3] ), .D(\Col_Fill[7][3] ), .S0(n65527), .S1(n65951), .Q(
        n3794) );
  IMUX21 U7273 ( .A(n3793), .B(n3794), .S(n65946), .Q(N1467) );
  IMUX40 U7499 ( .A(\Col_Fill[0][2] ), .B(\Col_Fill[1][2] ), .C(
        \Col_Fill[2][2] ), .D(\Col_Fill[3][2] ), .S0(n65516), .S1(n65940), .Q(
        n3919) );
  IMUX40 U7498 ( .A(\Col_Fill[4][2] ), .B(\Col_Fill[5][2] ), .C(
        \Col_Fill[6][2] ), .D(\Col_Fill[7][2] ), .S0(n65517), .S1(n65939), .Q(
        n3920) );
  IMUX21 U7464 ( .A(n3919), .B(n3920), .S(n65936), .Q(N2011) );
  IMUX40 U7307 ( .A(\Col_Fill[0][2] ), .B(\Col_Fill[1][2] ), .C(
        \Col_Fill[2][2] ), .D(\Col_Fill[3][2] ), .S0(n65529), .S1(n65950), .Q(
        n3791) );
  IMUX40 U7306 ( .A(\Col_Fill[4][2] ), .B(\Col_Fill[5][2] ), .C(
        \Col_Fill[6][2] ), .D(\Col_Fill[7][2] ), .S0(n65527), .S1(n65949), .Q(
        n3792) );
  IMUX21 U7272 ( .A(n3791), .B(n3792), .S(n65946), .Q(N1468) );
  IMUX40 U7497 ( .A(\Col_Fill[0][1] ), .B(\Col_Fill[1][1] ), .C(
        \Col_Fill[2][1] ), .D(\Col_Fill[3][1] ), .S0(n65419), .S1(n65943), .Q(
        n3917) );
  IMUX40 U7496 ( .A(\Col_Fill[4][1] ), .B(\Col_Fill[5][1] ), .C(
        \Col_Fill[6][1] ), .D(\Col_Fill[7][1] ), .S0(n65516), .S1(n65943), .Q(
        n3918) );
  IMUX21 U7463 ( .A(n3917), .B(n3918), .S(n65936), .Q(N2012) );
  IMUX40 U7305 ( .A(\Col_Fill[0][1] ), .B(\Col_Fill[1][1] ), .C(
        \Col_Fill[2][1] ), .D(\Col_Fill[3][1] ), .S0(n65525), .S1(n65953), .Q(
        n3789) );
  IMUX40 U7304 ( .A(\Col_Fill[4][1] ), .B(\Col_Fill[5][1] ), .C(
        \Col_Fill[6][1] ), .D(\Col_Fill[7][1] ), .S0(n65528), .S1(n65953), .Q(
        n3790) );
  IMUX21 U7271 ( .A(n3789), .B(n3790), .S(n65946), .Q(N1469) );
  IMUX40 U7555 ( .A(\Col_Fill[0][30] ), .B(\Col_Fill[1][30] ), .C(
        \Col_Fill[2][30] ), .D(\Col_Fill[3][30] ), .S0(n65518), .S1(n65940), 
        .Q(n3975) );
  IMUX40 U7554 ( .A(\Col_Fill[4][30] ), .B(\Col_Fill[5][30] ), .C(
        \Col_Fill[6][30] ), .D(\Col_Fill[7][30] ), .S0(n65521), .S1(n65938), 
        .Q(n3976) );
  IMUX21 U7492 ( .A(n3975), .B(n3976), .S(n65937), .Q(N1983) );
  IMUX40 U7363 ( .A(\Col_Fill[0][30] ), .B(\Col_Fill[1][30] ), .C(
        \Col_Fill[2][30] ), .D(\Col_Fill[3][30] ), .S0(n65531), .S1(n65950), 
        .Q(n3847) );
  IMUX40 U7362 ( .A(\Col_Fill[4][30] ), .B(\Col_Fill[5][30] ), .C(
        \Col_Fill[6][30] ), .D(\Col_Fill[7][30] ), .S0(n65531), .S1(n65948), 
        .Q(n3848) );
  IMUX21 U7300 ( .A(n3847), .B(n3848), .S(n65947), .Q(N1440) );
  IMUX40 U7557 ( .A(\Col_Fill[0][31] ), .B(\Col_Fill[1][31] ), .C(
        \Col_Fill[2][31] ), .D(\Col_Fill[3][31] ), .S0(n65419), .S1(n65938), 
        .Q(n3977) );
  IMUX40 U7556 ( .A(\Col_Fill[4][31] ), .B(\Col_Fill[5][31] ), .C(
        \Col_Fill[6][31] ), .D(\Col_Fill[7][31] ), .S0(n65520), .S1(n65939), 
        .Q(n3978) );
  IMUX21 U7493 ( .A(n3977), .B(n3978), .S(n65937), .Q(N1982) );
  IMUX40 U7365 ( .A(\Col_Fill[0][31] ), .B(\Col_Fill[1][31] ), .C(
        \Col_Fill[2][31] ), .D(\Col_Fill[3][31] ), .S0(n65531), .S1(n65948), 
        .Q(n3849) );
  IMUX40 U7364 ( .A(\Col_Fill[4][31] ), .B(\Col_Fill[5][31] ), .C(
        \Col_Fill[6][31] ), .D(\Col_Fill[7][31] ), .S0(n65531), .S1(n65949), 
        .Q(n3850) );
  IMUX21 U7301 ( .A(n3849), .B(n3850), .S(n65947), .Q(N1439) );
  IMUX40 U7207 ( .A(\Col_Fill[0][0] ), .B(\Col_Fill[1][0] ), .C(
        \Col_Fill[2][0] ), .D(\Col_Fill[3][0] ), .S0(n65527), .S1(n65953), .Q(
        n3723) );
  IMUX40 U7206 ( .A(\Col_Fill[4][0] ), .B(\Col_Fill[5][0] ), .C(
        \Col_Fill[6][0] ), .D(\Col_Fill[7][0] ), .S0(n65528), .S1(n65953), .Q(
        n3724) );
  IMUX21 U7174 ( .A(n3723), .B(n3724), .S(n65946), .Q(N1300) );
  IMUX40 U7399 ( .A(\Col_Fill[0][0] ), .B(\Col_Fill[1][0] ), .C(
        \Col_Fill[2][0] ), .D(\Col_Fill[3][0] ), .S0(n65517), .S1(n65943), .Q(
        n3851) );
  IMUX40 U7398 ( .A(\Col_Fill[4][0] ), .B(\Col_Fill[5][0] ), .C(
        \Col_Fill[6][0] ), .D(\Col_Fill[7][0] ), .S0(n65516), .S1(n65943), .Q(
        n3852) );
  IMUX21 U7366 ( .A(n3851), .B(n3852), .S(n65936), .Q(N1843) );
  IMUX40 U7495 ( .A(\Col_Fill[0][0] ), .B(\Col_Fill[1][0] ), .C(
        \Col_Fill[2][0] ), .D(\Col_Fill[3][0] ), .S0(n65517), .S1(n65943), .Q(
        n3915) );
  IMUX40 U7494 ( .A(\Col_Fill[4][0] ), .B(\Col_Fill[5][0] ), .C(
        \Col_Fill[6][0] ), .D(\Col_Fill[7][0] ), .S0(n65419), .S1(n65943), .Q(
        n3916) );
  IMUX21 U7462 ( .A(n3915), .B(n3916), .S(n65936), .Q(N2013) );
  IMUX40 U7303 ( .A(\Col_Fill[0][0] ), .B(\Col_Fill[1][0] ), .C(
        \Col_Fill[2][0] ), .D(\Col_Fill[3][0] ), .S0(n65527), .S1(n65953), .Q(
        n3787) );
  IMUX40 U7302 ( .A(\Col_Fill[4][0] ), .B(\Col_Fill[5][0] ), .C(
        \Col_Fill[6][0] ), .D(\Col_Fill[7][0] ), .S0(n65524), .S1(n65953), .Q(
        n3788) );
  IMUX21 U7270 ( .A(n3787), .B(n3788), .S(n65946), .Q(N1470) );
  IMUX40 U7411 ( .A(\Col_Fill[0][6] ), .B(\Col_Fill[1][6] ), .C(
        \Col_Fill[2][6] ), .D(\Col_Fill[3][6] ), .S0(n65516), .S1(n65940), .Q(
        n3863) );
  IMUX40 U7410 ( .A(\Col_Fill[4][6] ), .B(\Col_Fill[5][6] ), .C(
        \Col_Fill[6][6] ), .D(\Col_Fill[7][6] ), .S0(n65513), .S1(n65938), .Q(
        n3864) );
  IMUX21 U7372 ( .A(n3863), .B(n3864), .S(n65936), .Q(N1900) );
  IMUX40 U7219 ( .A(\Col_Fill[0][6] ), .B(\Col_Fill[1][6] ), .C(
        \Col_Fill[2][6] ), .D(\Col_Fill[3][6] ), .S0(n65526), .S1(n65950), .Q(
        n3735) );
  IMUX40 U7218 ( .A(\Col_Fill[4][6] ), .B(\Col_Fill[5][6] ), .C(
        \Col_Fill[6][6] ), .D(\Col_Fill[7][6] ), .S0(n65453), .S1(n65948), .Q(
        n3736) );
  IMUX21 U7180 ( .A(n3735), .B(n3736), .S(n65946), .Q(N1357) );
  IMUX40 U7441 ( .A(\Col_Fill[0][21] ), .B(\Col_Fill[1][21] ), .C(
        \Col_Fill[2][21] ), .D(\Col_Fill[3][21] ), .S0(n65512), .S1(n65944), 
        .Q(n3893) );
  IMUX40 U7440 ( .A(\Col_Fill[4][21] ), .B(\Col_Fill[5][21] ), .C(
        \Col_Fill[6][21] ), .D(\Col_Fill[7][21] ), .S0(n65511), .S1(n65945), 
        .Q(n3894) );
  IMUX21 U7387 ( .A(n3893), .B(n3894), .S(n65936), .Q(N1885) );
  IMUX40 U7249 ( .A(\Col_Fill[0][21] ), .B(\Col_Fill[1][21] ), .C(
        \Col_Fill[2][21] ), .D(\Col_Fill[3][21] ), .S0(n65526), .S1(n65954), 
        .Q(n3765) );
  IMUX40 U7248 ( .A(\Col_Fill[4][21] ), .B(\Col_Fill[5][21] ), .C(
        \Col_Fill[6][21] ), .D(\Col_Fill[7][21] ), .S0(n65524), .S1(n65955), 
        .Q(n3766) );
  IMUX21 U7195 ( .A(n3765), .B(n3766), .S(n65946), .Q(N1342) );
  IMUX40 U7221 ( .A(\Col_Fill[0][7] ), .B(\Col_Fill[1][7] ), .C(
        \Col_Fill[2][7] ), .D(\Col_Fill[3][7] ), .S0(n65527), .S1(n65951), .Q(
        n3737) );
  IMUX40 U7220 ( .A(\Col_Fill[4][7] ), .B(\Col_Fill[5][7] ), .C(
        \Col_Fill[6][7] ), .D(\Col_Fill[7][7] ), .S0(n65453), .S1(n65949), .Q(
        n3738) );
  IMUX21 U7181 ( .A(n3737), .B(n3738), .S(n65946), .Q(N1356) );
  IMUX40 U7413 ( .A(\Col_Fill[0][7] ), .B(\Col_Fill[1][7] ), .C(
        \Col_Fill[2][7] ), .D(\Col_Fill[3][7] ), .S0(n65522), .S1(n65941), .Q(
        n3865) );
  IMUX40 U7412 ( .A(\Col_Fill[4][7] ), .B(\Col_Fill[5][7] ), .C(
        \Col_Fill[6][7] ), .D(\Col_Fill[7][7] ), .S0(n65522), .S1(n65939), .Q(
        n3866) );
  IMUX21 U7373 ( .A(n3865), .B(n3866), .S(n65936), .Q(N1899) );
  IMUX40 U7267 ( .A(\Col_Fill[0][30] ), .B(\Col_Fill[1][30] ), .C(
        \Col_Fill[2][30] ), .D(\Col_Fill[3][30] ), .S0(n65530), .S1(n65955), 
        .Q(n3783) );
  IMUX40 U7266 ( .A(\Col_Fill[4][30] ), .B(\Col_Fill[5][30] ), .C(
        \Col_Fill[6][30] ), .D(\Col_Fill[7][30] ), .S0(n65453), .S1(n65955), 
        .Q(n3784) );
  IMUX21 U7204 ( .A(n3783), .B(n3784), .S(n65946), .Q(N1333) );
  IMUX40 U7459 ( .A(\Col_Fill[0][30] ), .B(\Col_Fill[1][30] ), .C(
        \Col_Fill[2][30] ), .D(\Col_Fill[3][30] ), .S0(n65510), .S1(n65945), 
        .Q(n3911) );
  IMUX40 U7458 ( .A(\Col_Fill[4][30] ), .B(\Col_Fill[5][30] ), .C(
        \Col_Fill[6][30] ), .D(\Col_Fill[7][30] ), .S0(n65515), .S1(n65945), 
        .Q(n3912) );
  IMUX21 U7396 ( .A(n3911), .B(n3912), .S(n65936), .Q(N1876) );
  IMUX40 U7217 ( .A(\Col_Fill[0][5] ), .B(\Col_Fill[1][5] ), .C(
        \Col_Fill[2][5] ), .D(\Col_Fill[3][5] ), .S0(n65532), .S1(n65950), .Q(
        n3733) );
  IMUX40 U7216 ( .A(\Col_Fill[4][5] ), .B(\Col_Fill[5][5] ), .C(
        \Col_Fill[6][5] ), .D(\Col_Fill[7][5] ), .S0(n65526), .S1(n65948), .Q(
        n3734) );
  IMUX21 U7179 ( .A(n3733), .B(n3734), .S(n65946), .Q(N1358) );
  IMUX40 U7437 ( .A(\Col_Fill[0][19] ), .B(\Col_Fill[1][19] ), .C(
        \Col_Fill[2][19] ), .D(\Col_Fill[3][19] ), .S0(n65511), .S1(n65943), 
        .Q(n3889) );
  IMUX40 U7436 ( .A(\Col_Fill[4][19] ), .B(\Col_Fill[5][19] ), .C(
        \Col_Fill[6][19] ), .D(\Col_Fill[7][19] ), .S0(n65516), .S1(n65942), 
        .Q(n3890) );
  IMUX21 U7385 ( .A(n3889), .B(n3890), .S(n65936), .Q(N1887) );
  IMUX40 U7409 ( .A(\Col_Fill[0][5] ), .B(\Col_Fill[1][5] ), .C(
        \Col_Fill[2][5] ), .D(\Col_Fill[3][5] ), .S0(n65515), .S1(n65940), .Q(
        n3861) );
  IMUX40 U7408 ( .A(\Col_Fill[4][5] ), .B(\Col_Fill[5][5] ), .C(
        \Col_Fill[6][5] ), .D(\Col_Fill[7][5] ), .S0(n65518), .S1(n65938), .Q(
        n3862) );
  IMUX21 U7371 ( .A(n3861), .B(n3862), .S(n65936), .Q(N1901) );
  IMUX40 U7245 ( .A(\Col_Fill[0][19] ), .B(\Col_Fill[1][19] ), .C(
        \Col_Fill[2][19] ), .D(\Col_Fill[3][19] ), .S0(n65524), .S1(n65953), 
        .Q(n3761) );
  IMUX40 U7244 ( .A(\Col_Fill[4][19] ), .B(\Col_Fill[5][19] ), .C(
        \Col_Fill[6][19] ), .D(\Col_Fill[7][19] ), .S0(n65527), .S1(n65952), 
        .Q(n3762) );
  IMUX21 U7193 ( .A(n3761), .B(n3762), .S(n65946), .Q(N1344) );
  IMUX40 U7239 ( .A(\Col_Fill[0][16] ), .B(\Col_Fill[1][16] ), .C(
        \Col_Fill[2][16] ), .D(\Col_Fill[3][16] ), .S0(n65420), .S1(n65948), 
        .Q(n3755) );
  IMUX40 U7238 ( .A(\Col_Fill[4][16] ), .B(\Col_Fill[5][16] ), .C(
        \Col_Fill[6][16] ), .D(\Col_Fill[7][16] ), .S0(n65525), .S1(n65951), 
        .Q(n3756) );
  IMUX21 U7190 ( .A(n3755), .B(n3756), .S(n65946), .Q(N1347) );
  IMUX40 U7431 ( .A(\Col_Fill[0][16] ), .B(\Col_Fill[1][16] ), .C(
        \Col_Fill[2][16] ), .D(\Col_Fill[3][16] ), .S0(n65419), .S1(n65938), 
        .Q(n3883) );
  IMUX40 U7430 ( .A(\Col_Fill[4][16] ), .B(\Col_Fill[5][16] ), .C(
        \Col_Fill[6][16] ), .D(\Col_Fill[7][16] ), .S0(n65516), .S1(n65941), 
        .Q(n3884) );
  IMUX21 U7382 ( .A(n3883), .B(n3884), .S(n65936), .Q(N1890) );
  IMUX40 U7415 ( .A(\Col_Fill[0][8] ), .B(\Col_Fill[1][8] ), .C(
        \Col_Fill[2][8] ), .D(\Col_Fill[3][8] ), .S0(n65515), .S1(N689), .Q(
        n3867) );
  IMUX40 U7414 ( .A(\Col_Fill[4][8] ), .B(\Col_Fill[5][8] ), .C(
        \Col_Fill[6][8] ), .D(\Col_Fill[7][8] ), .S0(n65514), .S1(n65939), .Q(
        n3868) );
  IMUX21 U7374 ( .A(n3867), .B(n3868), .S(n65936), .Q(N1898) );
  IMUX40 U7223 ( .A(\Col_Fill[0][8] ), .B(\Col_Fill[1][8] ), .C(
        \Col_Fill[2][8] ), .D(\Col_Fill[3][8] ), .S0(n65531), .S1(N683), .Q(
        n3739) );
  IMUX40 U7222 ( .A(\Col_Fill[4][8] ), .B(\Col_Fill[5][8] ), .C(
        \Col_Fill[6][8] ), .D(\Col_Fill[7][8] ), .S0(n65525), .S1(n65949), .Q(
        n3740) );
  IMUX21 U7182 ( .A(n3739), .B(n3740), .S(n65946), .Q(N1355) );
  IMUX40 U7439 ( .A(\Col_Fill[0][20] ), .B(\Col_Fill[1][20] ), .C(
        \Col_Fill[2][20] ), .D(\Col_Fill[3][20] ), .S0(n65513), .S1(n65940), 
        .Q(n3891) );
  IMUX40 U7438 ( .A(\Col_Fill[4][20] ), .B(\Col_Fill[5][20] ), .C(
        \Col_Fill[6][20] ), .D(\Col_Fill[7][20] ), .S0(n65512), .S1(n65939), 
        .Q(n3892) );
  IMUX21 U7386 ( .A(n3891), .B(n3892), .S(n65936), .Q(N1886) );
  IMUX40 U7247 ( .A(\Col_Fill[0][20] ), .B(\Col_Fill[1][20] ), .C(
        \Col_Fill[2][20] ), .D(\Col_Fill[3][20] ), .S0(n65527), .S1(n65950), 
        .Q(n3763) );
  IMUX40 U7246 ( .A(\Col_Fill[4][20] ), .B(\Col_Fill[5][20] ), .C(
        \Col_Fill[6][20] ), .D(\Col_Fill[7][20] ), .S0(n65530), .S1(n65949), 
        .Q(n3764) );
  IMUX21 U7194 ( .A(n3763), .B(n3764), .S(n65946), .Q(N1343) );
  IMUX40 U7263 ( .A(\Col_Fill[0][28] ), .B(\Col_Fill[1][28] ), .C(
        \Col_Fill[2][28] ), .D(\Col_Fill[3][28] ), .S0(n65530), .S1(n65955), 
        .Q(n3779) );
  IMUX40 U7262 ( .A(\Col_Fill[4][28] ), .B(\Col_Fill[5][28] ), .C(
        \Col_Fill[6][28] ), .D(\Col_Fill[7][28] ), .S0(n65523), .S1(n65955), 
        .Q(n3780) );
  IMUX21 U7202 ( .A(n3779), .B(n3780), .S(n65946), .Q(N1335) );
  IMUX40 U7455 ( .A(\Col_Fill[0][28] ), .B(\Col_Fill[1][28] ), .C(
        \Col_Fill[2][28] ), .D(\Col_Fill[3][28] ), .S0(n65517), .S1(n65945), 
        .Q(n3907) );
  IMUX40 U7454 ( .A(\Col_Fill[4][28] ), .B(\Col_Fill[5][28] ), .C(
        \Col_Fill[6][28] ), .D(\Col_Fill[7][28] ), .S0(n65512), .S1(n65945), 
        .Q(n3908) );
  IMUX21 U7394 ( .A(n3907), .B(n3908), .S(n65936), .Q(N1878) );
  IMUX40 U7231 ( .A(\Col_Fill[0][12] ), .B(\Col_Fill[1][12] ), .C(
        \Col_Fill[2][12] ), .D(\Col_Fill[3][12] ), .S0(n65525), .S1(n65954), 
        .Q(n3747) );
  IMUX40 U7230 ( .A(\Col_Fill[4][12] ), .B(\Col_Fill[5][12] ), .C(
        \Col_Fill[6][12] ), .D(\Col_Fill[7][12] ), .S0(n65525), .S1(n65954), 
        .Q(n3748) );
  IMUX21 U7186 ( .A(n3747), .B(n3748), .S(n65946), .Q(N1351) );
  IMUX40 U7423 ( .A(\Col_Fill[0][12] ), .B(\Col_Fill[1][12] ), .C(
        \Col_Fill[2][12] ), .D(\Col_Fill[3][12] ), .S0(n65514), .S1(n65944), 
        .Q(n3875) );
  IMUX40 U7422 ( .A(\Col_Fill[4][12] ), .B(\Col_Fill[5][12] ), .C(
        \Col_Fill[6][12] ), .D(\Col_Fill[7][12] ), .S0(n65515), .S1(n65944), 
        .Q(n3876) );
  IMUX21 U7378 ( .A(n3875), .B(n3876), .S(n65936), .Q(N1894) );
  IMUX40 U7241 ( .A(\Col_Fill[0][17] ), .B(\Col_Fill[1][17] ), .C(
        \Col_Fill[2][17] ), .D(\Col_Fill[3][17] ), .S0(n65453), .S1(n65954), 
        .Q(n3757) );
  IMUX40 U7240 ( .A(\Col_Fill[4][17] ), .B(\Col_Fill[5][17] ), .C(
        \Col_Fill[6][17] ), .D(\Col_Fill[7][17] ), .S0(n65525), .S1(n65955), 
        .Q(n3758) );
  IMUX21 U7191 ( .A(n3757), .B(n3758), .S(n65946), .Q(N1346) );
  IMUX40 U7269 ( .A(\Col_Fill[0][31] ), .B(\Col_Fill[1][31] ), .C(
        \Col_Fill[2][31] ), .D(\Col_Fill[3][31] ), .S0(n65527), .S1(n65955), 
        .Q(n3785) );
  IMUX40 U7268 ( .A(\Col_Fill[4][31] ), .B(\Col_Fill[5][31] ), .C(
        \Col_Fill[6][31] ), .D(\Col_Fill[7][31] ), .S0(n65523), .S1(n65955), 
        .Q(n3786) );
  IMUX21 U7205 ( .A(n3785), .B(n3786), .S(n65946), .Q(N1332) );
  IMUX40 U7225 ( .A(\Col_Fill[0][9] ), .B(\Col_Fill[1][9] ), .C(
        \Col_Fill[2][9] ), .D(\Col_Fill[3][9] ), .S0(n65525), .S1(n65948), .Q(
        n3741) );
  IMUX40 U7224 ( .A(\Col_Fill[4][9] ), .B(\Col_Fill[5][9] ), .C(
        \Col_Fill[6][9] ), .D(\Col_Fill[7][9] ), .S0(n65523), .S1(n65951), .Q(
        n3742) );
  IMUX21 U7183 ( .A(n3741), .B(n3742), .S(n65946), .Q(N1354) );
  IMUX40 U7417 ( .A(\Col_Fill[0][9] ), .B(\Col_Fill[1][9] ), .C(
        \Col_Fill[2][9] ), .D(\Col_Fill[3][9] ), .S0(n65514), .S1(n65938), .Q(
        n3869) );
  IMUX40 U7416 ( .A(\Col_Fill[4][9] ), .B(\Col_Fill[5][9] ), .C(
        \Col_Fill[6][9] ), .D(\Col_Fill[7][9] ), .S0(n65517), .S1(n65941), .Q(
        n3870) );
  IMUX21 U7375 ( .A(n3869), .B(n3870), .S(n65936), .Q(N1897) );
  IMUX40 U7259 ( .A(\Col_Fill[0][26] ), .B(\Col_Fill[1][26] ), .C(
        \Col_Fill[2][26] ), .D(\Col_Fill[3][26] ), .S0(n65523), .S1(n65951), 
        .Q(n3775) );
  IMUX40 U7258 ( .A(\Col_Fill[4][26] ), .B(\Col_Fill[5][26] ), .C(
        \Col_Fill[6][26] ), .D(\Col_Fill[7][26] ), .S0(n65420), .S1(N683), .Q(
        n3776) );
  IMUX21 U7200 ( .A(n3775), .B(n3776), .S(n65946), .Q(N1337) );
  IMUX40 U7461 ( .A(\Col_Fill[0][31] ), .B(\Col_Fill[1][31] ), .C(
        \Col_Fill[2][31] ), .D(\Col_Fill[3][31] ), .S0(n65517), .S1(n65945), 
        .Q(n3913) );
  IMUX40 U7460 ( .A(\Col_Fill[4][31] ), .B(\Col_Fill[5][31] ), .C(
        \Col_Fill[6][31] ), .D(\Col_Fill[7][31] ), .S0(n65519), .S1(n65945), 
        .Q(n3914) );
  IMUX21 U7397 ( .A(n3913), .B(n3914), .S(n65936), .Q(N1875) );
  IMUX40 U7451 ( .A(\Col_Fill[0][26] ), .B(\Col_Fill[1][26] ), .C(
        \Col_Fill[2][26] ), .D(\Col_Fill[3][26] ), .S0(n65520), .S1(n65941), 
        .Q(n3903) );
  IMUX40 U7450 ( .A(\Col_Fill[4][26] ), .B(\Col_Fill[5][26] ), .C(
        \Col_Fill[6][26] ), .D(\Col_Fill[7][26] ), .S0(n65510), .S1(N689), .Q(
        n3904) );
  IMUX21 U7392 ( .A(n3903), .B(n3904), .S(n65936), .Q(N1880) );
  IMUX40 U7433 ( .A(\Col_Fill[0][17] ), .B(\Col_Fill[1][17] ), .C(
        \Col_Fill[2][17] ), .D(\Col_Fill[3][17] ), .S0(n65516), .S1(n65944), 
        .Q(n3885) );
  IMUX40 U7432 ( .A(\Col_Fill[4][17] ), .B(\Col_Fill[5][17] ), .C(
        \Col_Fill[6][17] ), .D(\Col_Fill[7][17] ), .S0(n65419), .S1(n65945), 
        .Q(n3886) );
  IMUX21 U7383 ( .A(n3885), .B(n3886), .S(n65936), .Q(N1889) );
  IMUX40 U7445 ( .A(\Col_Fill[0][23] ), .B(\Col_Fill[1][23] ), .C(
        \Col_Fill[2][23] ), .D(\Col_Fill[3][23] ), .S0(n65513), .S1(n65938), 
        .Q(n3897) );
  IMUX40 U7444 ( .A(\Col_Fill[4][23] ), .B(\Col_Fill[5][23] ), .C(
        \Col_Fill[6][23] ), .D(\Col_Fill[7][23] ), .S0(n65512), .S1(n65940), 
        .Q(n3898) );
  IMUX21 U7389 ( .A(n3897), .B(n3898), .S(n65936), .Q(N1883) );
  IMUX40 U7253 ( .A(\Col_Fill[0][23] ), .B(\Col_Fill[1][23] ), .C(
        \Col_Fill[2][23] ), .D(\Col_Fill[3][23] ), .S0(n65531), .S1(n65948), 
        .Q(n3769) );
  IMUX40 U7252 ( .A(\Col_Fill[4][23] ), .B(\Col_Fill[5][23] ), .C(
        \Col_Fill[6][23] ), .D(\Col_Fill[7][23] ), .S0(n65529), .S1(n65950), 
        .Q(n3770) );
  IMUX21 U7197 ( .A(n3769), .B(n3770), .S(n65946), .Q(N1340) );
  IMUX40 U7265 ( .A(\Col_Fill[0][29] ), .B(\Col_Fill[1][29] ), .C(
        \Col_Fill[2][29] ), .D(\Col_Fill[3][29] ), .S0(n65523), .S1(n65955), 
        .Q(n3781) );
  IMUX40 U7264 ( .A(\Col_Fill[4][29] ), .B(\Col_Fill[5][29] ), .C(
        \Col_Fill[6][29] ), .D(\Col_Fill[7][29] ), .S0(n65524), .S1(n65955), 
        .Q(n3782) );
  IMUX21 U7203 ( .A(n3781), .B(n3782), .S(n65946), .Q(N1334) );
  IMUX40 U7457 ( .A(\Col_Fill[0][29] ), .B(\Col_Fill[1][29] ), .C(
        \Col_Fill[2][29] ), .D(\Col_Fill[3][29] ), .S0(n65519), .S1(n65945), 
        .Q(n3909) );
  IMUX40 U7456 ( .A(\Col_Fill[4][29] ), .B(\Col_Fill[5][29] ), .C(
        \Col_Fill[6][29] ), .D(\Col_Fill[7][29] ), .S0(n65510), .S1(n65945), 
        .Q(n3910) );
  IMUX21 U7395 ( .A(n3909), .B(n3910), .S(n65936), .Q(N1877) );
  IMUX40 U7237 ( .A(\Col_Fill[0][15] ), .B(\Col_Fill[1][15] ), .C(
        \Col_Fill[2][15] ), .D(\Col_Fill[3][15] ), .S0(n65531), .S1(n65954), 
        .Q(n3753) );
  IMUX40 U7236 ( .A(\Col_Fill[4][15] ), .B(\Col_Fill[5][15] ), .C(
        \Col_Fill[6][15] ), .D(\Col_Fill[7][15] ), .S0(n65420), .S1(n65954), 
        .Q(n3754) );
  IMUX21 U7189 ( .A(n3753), .B(n3754), .S(n65946), .Q(N1348) );
  IMUX40 U7429 ( .A(\Col_Fill[0][15] ), .B(\Col_Fill[1][15] ), .C(
        \Col_Fill[2][15] ), .D(\Col_Fill[3][15] ), .S0(n65517), .S1(n65944), 
        .Q(n3881) );
  IMUX40 U7428 ( .A(\Col_Fill[4][15] ), .B(\Col_Fill[5][15] ), .C(
        \Col_Fill[6][15] ), .D(\Col_Fill[7][15] ), .S0(n65518), .S1(n65944), 
        .Q(n3882) );
  IMUX21 U7381 ( .A(n3881), .B(n3882), .S(n65936), .Q(N1891) );
  IMUX40 U7235 ( .A(\Col_Fill[0][14] ), .B(\Col_Fill[1][14] ), .C(
        \Col_Fill[2][14] ), .D(\Col_Fill[3][14] ), .S0(n65529), .S1(n65954), 
        .Q(n3751) );
  IMUX40 U7234 ( .A(\Col_Fill[4][14] ), .B(\Col_Fill[5][14] ), .C(
        \Col_Fill[6][14] ), .D(\Col_Fill[7][14] ), .S0(n65523), .S1(n65954), 
        .Q(n3752) );
  IMUX21 U7188 ( .A(n3751), .B(n3752), .S(n65946), .Q(N1349) );
  IMUX40 U7427 ( .A(\Col_Fill[0][14] ), .B(\Col_Fill[1][14] ), .C(
        \Col_Fill[2][14] ), .D(\Col_Fill[3][14] ), .S0(n65419), .S1(n65944), 
        .Q(n3879) );
  IMUX40 U7426 ( .A(\Col_Fill[4][14] ), .B(\Col_Fill[5][14] ), .C(
        \Col_Fill[6][14] ), .D(\Col_Fill[7][14] ), .S0(n65511), .S1(n65944), 
        .Q(n3880) );
  IMUX21 U7380 ( .A(n3879), .B(n3880), .S(n65936), .Q(N1892) );
  IMUX40 U7233 ( .A(\Col_Fill[0][13] ), .B(\Col_Fill[1][13] ), .C(
        \Col_Fill[2][13] ), .D(\Col_Fill[3][13] ), .S0(n65420), .S1(n65954), 
        .Q(n3749) );
  IMUX40 U7232 ( .A(\Col_Fill[4][13] ), .B(\Col_Fill[5][13] ), .C(
        \Col_Fill[6][13] ), .D(\Col_Fill[7][13] ), .S0(n65526), .S1(n65954), 
        .Q(n3750) );
  IMUX21 U7187 ( .A(n3749), .B(n3750), .S(n65946), .Q(N1350) );
  IMUX40 U7425 ( .A(\Col_Fill[0][13] ), .B(\Col_Fill[1][13] ), .C(
        \Col_Fill[2][13] ), .D(\Col_Fill[3][13] ), .S0(n65521), .S1(n65944), 
        .Q(n3877) );
  IMUX40 U7424 ( .A(\Col_Fill[4][13] ), .B(\Col_Fill[5][13] ), .C(
        \Col_Fill[6][13] ), .D(\Col_Fill[7][13] ), .S0(n65515), .S1(n65944), 
        .Q(n3878) );
  IMUX21 U7379 ( .A(n3877), .B(n3878), .S(n65936), .Q(N1893) );
  IMUX40 U7261 ( .A(\Col_Fill[0][27] ), .B(\Col_Fill[1][27] ), .C(
        \Col_Fill[2][27] ), .D(\Col_Fill[3][27] ), .S0(n65453), .S1(N683), .Q(
        n3777) );
  IMUX40 U7260 ( .A(\Col_Fill[4][27] ), .B(\Col_Fill[5][27] ), .C(
        \Col_Fill[6][27] ), .D(\Col_Fill[7][27] ), .S0(n65528), .S1(n65949), 
        .Q(n3778) );
  IMUX21 U7201 ( .A(n3777), .B(n3778), .S(n65946), .Q(N1336) );
  IMUX40 U7453 ( .A(\Col_Fill[0][27] ), .B(\Col_Fill[1][27] ), .C(
        \Col_Fill[2][27] ), .D(\Col_Fill[3][27] ), .S0(n65510), .S1(N689), .Q(
        n3905) );
  IMUX40 U7452 ( .A(\Col_Fill[4][27] ), .B(\Col_Fill[5][27] ), .C(
        \Col_Fill[6][27] ), .D(\Col_Fill[7][27] ), .S0(n65513), .S1(n65939), 
        .Q(n3906) );
  IMUX21 U7393 ( .A(n3905), .B(n3906), .S(n65936), .Q(N1879) );
  IMUX40 U7435 ( .A(\Col_Fill[0][18] ), .B(\Col_Fill[1][18] ), .C(
        \Col_Fill[2][18] ), .D(\Col_Fill[3][18] ), .S0(n65513), .S1(n65943), 
        .Q(n3887) );
  IMUX40 U7434 ( .A(\Col_Fill[4][18] ), .B(\Col_Fill[5][18] ), .C(
        \Col_Fill[6][18] ), .D(\Col_Fill[7][18] ), .S0(n65510), .S1(n65942), 
        .Q(n3888) );
  IMUX21 U7384 ( .A(n3887), .B(n3888), .S(n65936), .Q(N1888) );
  IMUX40 U7243 ( .A(\Col_Fill[0][18] ), .B(\Col_Fill[1][18] ), .C(
        \Col_Fill[2][18] ), .D(\Col_Fill[3][18] ), .S0(n65532), .S1(n65953), 
        .Q(n3759) );
  IMUX40 U7242 ( .A(\Col_Fill[4][18] ), .B(\Col_Fill[5][18] ), .C(
        \Col_Fill[6][18] ), .D(\Col_Fill[7][18] ), .S0(n65420), .S1(n65952), 
        .Q(n3760) );
  IMUX21 U7192 ( .A(n3759), .B(n3760), .S(n65946), .Q(N1345) );
  IMUX40 U7443 ( .A(\Col_Fill[0][22] ), .B(\Col_Fill[1][22] ), .C(
        \Col_Fill[2][22] ), .D(\Col_Fill[3][22] ), .S0(n65511), .S1(n65940), 
        .Q(n3895) );
  IMUX40 U7442 ( .A(\Col_Fill[4][22] ), .B(\Col_Fill[5][22] ), .C(
        \Col_Fill[6][22] ), .D(\Col_Fill[7][22] ), .S0(n65513), .S1(n65941), 
        .Q(n3896) );
  IMUX21 U7388 ( .A(n3895), .B(n3896), .S(n65936), .Q(N1884) );
  IMUX40 U7251 ( .A(\Col_Fill[0][22] ), .B(\Col_Fill[1][22] ), .C(
        \Col_Fill[2][22] ), .D(\Col_Fill[3][22] ), .S0(n65524), .S1(n65950), 
        .Q(n3767) );
  IMUX40 U7250 ( .A(\Col_Fill[4][22] ), .B(\Col_Fill[5][22] ), .C(
        \Col_Fill[6][22] ), .D(\Col_Fill[7][22] ), .S0(n65523), .S1(n65951), 
        .Q(n3768) );
  IMUX21 U7196 ( .A(n3767), .B(n3768), .S(n65946), .Q(N1341) );
  IMUX40 U7257 ( .A(\Col_Fill[0][25] ), .B(\Col_Fill[1][25] ), .C(
        \Col_Fill[2][25] ), .D(\Col_Fill[3][25] ), .S0(n65533), .S1(n65949), 
        .Q(n3773) );
  IMUX40 U7256 ( .A(\Col_Fill[4][25] ), .B(\Col_Fill[5][25] ), .C(
        \Col_Fill[6][25] ), .D(\Col_Fill[7][25] ), .S0(n65420), .S1(n65948), 
        .Q(n3774) );
  IMUX21 U7199 ( .A(n3773), .B(n3774), .S(n65946), .Q(N1338) );
  IMUX40 U7449 ( .A(\Col_Fill[0][25] ), .B(\Col_Fill[1][25] ), .C(
        \Col_Fill[2][25] ), .D(\Col_Fill[3][25] ), .S0(n65514), .S1(n65939), 
        .Q(n3901) );
  IMUX40 U7448 ( .A(\Col_Fill[4][25] ), .B(\Col_Fill[5][25] ), .C(
        \Col_Fill[6][25] ), .D(\Col_Fill[7][25] ), .S0(n65513), .S1(n65938), 
        .Q(n3902) );
  IMUX21 U7391 ( .A(n3901), .B(n3902), .S(n65936), .Q(N1881) );
  IMUX40 U7229 ( .A(\Col_Fill[0][11] ), .B(\Col_Fill[1][11] ), .C(
        \Col_Fill[2][11] ), .D(\Col_Fill[3][11] ), .S0(n65531), .S1(n65954), 
        .Q(n3745) );
  IMUX40 U7228 ( .A(\Col_Fill[4][11] ), .B(\Col_Fill[5][11] ), .C(
        \Col_Fill[6][11] ), .D(\Col_Fill[7][11] ), .S0(n65525), .S1(n65954), 
        .Q(n3746) );
  IMUX21 U7185 ( .A(n3745), .B(n3746), .S(n65946), .Q(N1352) );
  IMUX40 U7421 ( .A(\Col_Fill[0][11] ), .B(\Col_Fill[1][11] ), .C(
        \Col_Fill[2][11] ), .D(\Col_Fill[3][11] ), .S0(n65515), .S1(n65944), 
        .Q(n3873) );
  IMUX40 U7420 ( .A(\Col_Fill[4][11] ), .B(\Col_Fill[5][11] ), .C(
        \Col_Fill[6][11] ), .D(\Col_Fill[7][11] ), .S0(n65514), .S1(n65944), 
        .Q(n3874) );
  IMUX21 U7377 ( .A(n3873), .B(n3874), .S(n65936), .Q(N1895) );
  IMUX40 U7227 ( .A(\Col_Fill[0][10] ), .B(\Col_Fill[1][10] ), .C(
        \Col_Fill[2][10] ), .D(\Col_Fill[3][10] ), .S0(n65526), .S1(n65954), 
        .Q(n3743) );
  IMUX40 U7226 ( .A(\Col_Fill[4][10] ), .B(\Col_Fill[5][10] ), .C(
        \Col_Fill[6][10] ), .D(\Col_Fill[7][10] ), .S0(n65529), .S1(n65954), 
        .Q(n3744) );
  IMUX21 U7184 ( .A(n3743), .B(n3744), .S(n65946), .Q(N1353) );
  IMUX40 U7419 ( .A(\Col_Fill[0][10] ), .B(\Col_Fill[1][10] ), .C(
        \Col_Fill[2][10] ), .D(\Col_Fill[3][10] ), .S0(n65513), .S1(n65944), 
        .Q(n3871) );
  IMUX40 U7418 ( .A(\Col_Fill[4][10] ), .B(\Col_Fill[5][10] ), .C(
        \Col_Fill[6][10] ), .D(\Col_Fill[7][10] ), .S0(n65515), .S1(n65944), 
        .Q(n3872) );
  IMUX21 U7376 ( .A(n3871), .B(n3872), .S(n65936), .Q(N1896) );
  IMUX40 U7255 ( .A(\Col_Fill[0][24] ), .B(\Col_Fill[1][24] ), .C(
        \Col_Fill[2][24] ), .D(\Col_Fill[3][24] ), .S0(n65420), .S1(n65951), 
        .Q(n3771) );
  IMUX40 U7254 ( .A(\Col_Fill[4][24] ), .B(\Col_Fill[5][24] ), .C(
        \Col_Fill[6][24] ), .D(\Col_Fill[7][24] ), .S0(n65524), .S1(n65951), 
        .Q(n3772) );
  IMUX21 U7198 ( .A(n3771), .B(n3772), .S(n65946), .Q(N1339) );
  IMUX40 U7447 ( .A(\Col_Fill[0][24] ), .B(\Col_Fill[1][24] ), .C(
        \Col_Fill[2][24] ), .D(\Col_Fill[3][24] ), .S0(n65512), .S1(n65941), 
        .Q(n3899) );
  IMUX40 U7446 ( .A(\Col_Fill[4][24] ), .B(\Col_Fill[5][24] ), .C(
        \Col_Fill[6][24] ), .D(\Col_Fill[7][24] ), .S0(n65511), .S1(n65941), 
        .Q(n3900) );
  IMUX21 U7390 ( .A(n3899), .B(n3900), .S(n65936), .Q(N1882) );
  IMUX40 U7401 ( .A(\Col_Fill[0][1] ), .B(\Col_Fill[1][1] ), .C(
        \Col_Fill[2][1] ), .D(\Col_Fill[3][1] ), .S0(n65514), .S1(n65943), .Q(
        n3853) );
  IMUX40 U7400 ( .A(\Col_Fill[4][1] ), .B(\Col_Fill[5][1] ), .C(
        \Col_Fill[6][1] ), .D(\Col_Fill[7][1] ), .S0(n65510), .S1(n65943), .Q(
        n3854) );
  IMUX21 U7367 ( .A(n3853), .B(n3854), .S(n65936), .Q(N1905) );
  IMUX40 U7407 ( .A(\Col_Fill[0][4] ), .B(\Col_Fill[1][4] ), .C(
        \Col_Fill[2][4] ), .D(\Col_Fill[3][4] ), .S0(n65512), .S1(n65940), .Q(
        n3859) );
  IMUX40 U7406 ( .A(\Col_Fill[4][4] ), .B(\Col_Fill[5][4] ), .C(
        \Col_Fill[6][4] ), .D(\Col_Fill[7][4] ), .S0(n65517), .S1(n65940), .Q(
        n3860) );
  IMUX40 U7213 ( .A(\Col_Fill[0][3] ), .B(\Col_Fill[1][3] ), .C(
        \Col_Fill[2][3] ), .D(\Col_Fill[3][3] ), .S0(n65526), .S1(n65953), .Q(
        n3729) );
  IMUX40 U7212 ( .A(\Col_Fill[4][3] ), .B(\Col_Fill[5][3] ), .C(
        \Col_Fill[6][3] ), .D(\Col_Fill[7][3] ), .S0(n65529), .S1(n65953), .Q(
        n3730) );
  IMUX40 U7211 ( .A(\Col_Fill[0][2] ), .B(\Col_Fill[1][2] ), .C(
        \Col_Fill[2][2] ), .D(\Col_Fill[3][2] ), .S0(n65530), .S1(n65953), .Q(
        n3727) );
  IMUX40 U7210 ( .A(\Col_Fill[4][2] ), .B(\Col_Fill[5][2] ), .C(
        \Col_Fill[6][2] ), .D(\Col_Fill[7][2] ), .S0(n65526), .S1(n65953), .Q(
        n3728) );
  IMUX40 U7209 ( .A(\Col_Fill[0][1] ), .B(\Col_Fill[1][1] ), .C(
        \Col_Fill[2][1] ), .D(\Col_Fill[3][1] ), .S0(n65528), .S1(n65953), .Q(
        n3725) );
  IMUX40 U7208 ( .A(\Col_Fill[4][1] ), .B(\Col_Fill[5][1] ), .C(
        \Col_Fill[6][1] ), .D(\Col_Fill[7][1] ), .S0(n65523), .S1(n65953), .Q(
        n3726) );
  IMUX40 U7215 ( .A(\Col_Fill[0][4] ), .B(\Col_Fill[1][4] ), .C(
        \Col_Fill[2][4] ), .D(\Col_Fill[3][4] ), .S0(n65533), .S1(n65950), .Q(
        n3731) );
  IMUX40 U7214 ( .A(\Col_Fill[4][4] ), .B(\Col_Fill[5][4] ), .C(
        \Col_Fill[6][4] ), .D(\Col_Fill[7][4] ), .S0(n65523), .S1(n65950), .Q(
        n3732) );
  IMUX40 U7405 ( .A(\Col_Fill[0][3] ), .B(\Col_Fill[1][3] ), .C(
        \Col_Fill[2][3] ), .D(\Col_Fill[3][3] ), .S0(n65521), .S1(n65943), .Q(
        n3857) );
  IMUX40 U7404 ( .A(\Col_Fill[4][3] ), .B(\Col_Fill[5][3] ), .C(
        \Col_Fill[6][3] ), .D(\Col_Fill[7][3] ), .S0(n65519), .S1(n65943), .Q(
        n3858) );
  IMUX40 U7403 ( .A(\Col_Fill[0][2] ), .B(\Col_Fill[1][2] ), .C(
        \Col_Fill[2][2] ), .D(\Col_Fill[3][2] ), .S0(n65513), .S1(n65943), .Q(
        n3855) );
  IMUX40 U7402 ( .A(\Col_Fill[4][2] ), .B(\Col_Fill[5][2] ), .C(
        \Col_Fill[6][2] ), .D(\Col_Fill[7][2] ), .S0(n65510), .S1(n65943), .Q(
        n3856) );
  MUX41 U26378 ( .A(n21914), .B(n21904), .C(n21909), .D(n21899), .S0(N864), 
        .S1(N863), .Q(N4261) );
  MUX41 U58634 ( .A(n52634), .B(n52624), .C(n52629), .D(n52619), .S0(N1152), 
        .S1(N1151), .Q(N6531) );
  MUX41 U36458 ( .A(n31514), .B(n31504), .C(n31509), .D(n31499), .S0(N954), 
        .S1(N953), .Q(N4952) );
  MUX41 U68714 ( .A(n62234), .B(n62224), .C(n62229), .D(n62219), .S0(N1242), 
        .S1(N1241), .Q(N7222) );
  MUX41 U56618 ( .A(n50714), .B(n50704), .C(n50709), .D(n50699), .S0(N1134), 
        .S1(N1133), .Q(N6394) );
  IMUX40 U70054 ( .A(n63500), .B(n63501), .C(n63502), .D(n63503), .S0(N1252), 
        .S1(n65916), .Q(n63499) );
  IMUX40 U70055 ( .A(n63505), .B(n63506), .C(n63507), .D(n63508), .S0(N1252), 
        .S1(n65916), .Q(n63504) );
  MUX41 U70058 ( .A(n63514), .B(n63504), .C(n63509), .D(n63499), .S0(N1254), 
        .S1(N1253), .Q(N7328) );
  IMUX40 U37798 ( .A(n32780), .B(n32781), .C(n32782), .D(n32783), .S0(N964), 
        .S1(n65916), .Q(n32779) );
  IMUX40 U37799 ( .A(n32785), .B(n32786), .C(n32787), .D(n32788), .S0(N964), 
        .S1(n65916), .Q(n32784) );
  MUX41 U37802 ( .A(n32794), .B(n32784), .C(n32789), .D(n32779), .S0(N966), 
        .S1(N965), .Q(N5058) );
  IMUX40 U35110 ( .A(n30220), .B(n30221), .C(n30222), .D(n30223), .S0(N940), 
        .S1(n65918), .Q(n30219) );
  IMUX40 U35111 ( .A(n30225), .B(n30226), .C(n30227), .D(n30228), .S0(N940), 
        .S1(n65918), .Q(n30224) );
  MUX41 U35114 ( .A(n30234), .B(n30224), .C(n30229), .D(n30219), .S0(N942), 
        .S1(N941), .Q(N4845) );
  IMUX40 U67366 ( .A(n60940), .B(n60941), .C(n60942), .D(n60943), .S0(N1228), 
        .S1(n65917), .Q(n60939) );
  IMUX40 U67367 ( .A(n60945), .B(n60946), .C(n60947), .D(n60948), .S0(N1228), 
        .S1(n65917), .Q(n60944) );
  MUX41 U67370 ( .A(n60954), .B(n60944), .C(n60949), .D(n60939), .S0(N1230), 
        .S1(N1229), .Q(N7115) );
  MUX41 U39818 ( .A(n34714), .B(n34704), .C(n34709), .D(n34699), .S0(N984), 
        .S1(N983), .Q(N5246) );
  MUX41 U40490 ( .A(n35354), .B(n35344), .C(n35349), .D(n35339), .S0(N990), 
        .S1(N989), .Q(N5278) );
  MUX41 U25034 ( .A(n20634), .B(n20624), .C(n20629), .D(n20619), .S0(N852), 
        .S1(N851), .Q(N4156) );
  MUX41 U39146 ( .A(n34074), .B(n34064), .C(n34069), .D(n34059), .S0(N978), 
        .S1(N977), .Q(N5122) );
  MUX41 U12938 ( .A(n9114), .B(n9104), .C(n9109), .D(n9099), .S0(N744), .S1(
        N743), .Q(N3349) );
  MUX41 U64682 ( .A(n58394), .B(n58384), .C(n58389), .D(n58379), .S0(N1206), 
        .S1(N1205), .Q(N6946) );
  IMUX40 U37963 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65877), 
        .S1(n65753), .Q(n32786) );
  IMUX40 U37962 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65877), 
        .S1(n65745), .Q(n32788) );
  IMUX40 U37959 ( .A(n65684), .B(n65685), .C(n65686), .D(n65687), .S0(n65878), 
        .S1(n65752), .Q(n32781) );
  IMUX40 U37958 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(n65879), 
        .S1(n65755), .Q(n32783) );
  IMUX40 U35947 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65873), 
        .S1(n65762), .Q(n30866) );
  IMUX40 U35946 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65874), 
        .S1(n65763), .Q(n30868) );
  IMUX40 U35943 ( .A(n65684), .B(n65685), .C(n65686), .D(n65687), .S0(n65900), 
        .S1(n65778), .Q(n30861) );
  IMUX40 U35942 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(n65892), 
        .S1(n65770), .Q(n30863) );
  IMUX40 U35955 ( .A(n65732), .B(n65733), .C(n65734), .D(n65735), .S0(n65872), 
        .S1(n65780), .Q(n30876) );
  IMUX40 U35954 ( .A(n65736), .B(n65737), .C(n65738), .D(n65739), .S0(n65850), 
        .S1(n65771), .Q(n30878) );
  IMUX40 U70219 ( .A(n65636), .B(n65637), .C(n65638), .D(n65639), .S0(n65907), 
        .S1(n65753), .Q(n63506) );
  IMUX40 U70218 ( .A(n65640), .B(n65641), .C(n65642), .D(n65643), .S0(n65832), 
        .S1(n65753), .Q(n63508) );
  IMUX40 U70215 ( .A(n65620), .B(n65621), .C(n65622), .D(n65623), .S0(n65839), 
        .S1(n65753), .Q(n63501) );
  IMUX40 U70214 ( .A(n65624), .B(n65625), .C(n65626), .D(n65627), .S0(n65891), 
        .S1(n65753), .Q(n63503) );
  IMUX40 U71563 ( .A(n65636), .B(n65637), .C(n65638), .D(n65639), .S0(n65884), 
        .S1(n65765), .Q(n64786) );
  IMUX40 U71562 ( .A(n65640), .B(n65641), .C(n65642), .D(n65643), .S0(n65888), 
        .S1(n65765), .Q(n64788) );
  IMUX40 U71559 ( .A(n65620), .B(n65621), .C(n65622), .D(n65623), .S0(n65875), 
        .S1(n65765), .Q(n64781) );
  IMUX40 U71558 ( .A(n65624), .B(n65625), .C(n65626), .D(n65627), .S0(n65838), 
        .S1(n65764), .Q(n64783) );
  IMUX40 U68203 ( .A(n65636), .B(n65637), .C(n65638), .D(n65639), .S0(n65843), 
        .S1(n65768), .Q(n61586) );
  IMUX40 U68202 ( .A(n65640), .B(n65641), .C(n65642), .D(n65643), .S0(n65845), 
        .S1(n65767), .Q(n61588) );
  IMUX40 U68199 ( .A(n65620), .B(n65621), .C(n65622), .D(n65623), .S0(n65864), 
        .S1(n65772), .Q(n61581) );
  IMUX40 U68198 ( .A(n65624), .B(n65625), .C(n65626), .D(n65627), .S0(n65855), 
        .S1(n65780), .Q(n61583) );
  IMUX40 U68211 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65890), 
        .S1(n65759), .Q(n61596) );
  IMUX40 U68210 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65909), 
        .S1(n65773), .Q(n61598) );
  IMUX40 U70891 ( .A(n65636), .B(n65637), .C(n65638), .D(n65639), .S0(n65785), 
        .S1(N1256), .Q(n64146) );
  IMUX40 U70890 ( .A(n65640), .B(n65641), .C(n65642), .D(n65643), .S0(n65828), 
        .S1(N1256), .Q(n64148) );
  IMUX40 U70887 ( .A(n65620), .B(n65621), .C(n65622), .D(n65623), .S0(n65811), 
        .S1(N1256), .Q(n64141) );
  IMUX40 U70886 ( .A(n65624), .B(n65625), .C(n65626), .D(n65627), .S0(n65805), 
        .S1(N1256), .Q(n64143) );
  IMUX40 U70899 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65811), 
        .S1(N1256), .Q(n64156) );
  IMUX40 U70898 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65809), 
        .S1(N1256), .Q(n64158) );
  IMUX40 U49387 ( .A(\OFill[40][0] ), .B(n65637), .C(n65638), .D(n65639), .S0(
        n65894), .S1(n65749), .Q(n43666) );
  IMUX40 U49386 ( .A(\OFill[44][0] ), .B(n65641), .C(n65642), .D(n65643), .S0(
        n65889), .S1(n65751), .Q(n43668) );
  IMUX40 U49383 ( .A(\OFill[56][0] ), .B(n65621), .C(n65622), .D(n65623), .S0(
        n65897), .S1(n65749), .Q(n43661) );
  IMUX40 U49382 ( .A(\OFill[60][0] ), .B(n65625), .C(n65626), .D(n65627), .S0(
        n65896), .S1(n65754), .Q(n43663) );
  IMUX40 U49395 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65909), 
        .S1(n65750), .Q(n43676) );
  IMUX40 U49394 ( .A(n65672), .B(\OFill[13][0] ), .C(n65674), .D(n65675), .S0(
        n65900), .S1(n65756), .Q(n43678) );
  IMUX40 U50059 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65840), .S1(N1208), .Q(n44306) );
  IMUX40 U50058 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65840), .S1(n65748), .Q(n44308) );
  IMUX40 U50055 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65839), .S1(n65744), .Q(n44301) );
  IMUX40 U50054 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65839), .S1(n65746), .Q(n44303) );
  IMUX40 U50067 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65843), .S1(n65748), .Q(n44316) );
  IMUX40 U50066 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65843), .S1(n65757), .Q(n44318) );
  IMUX40 U51403 ( .A(n65636), .B(n65637), .C(n65638), .D(n65639), .S0(n65816), 
        .S1(n65912), .Q(n45586) );
  IMUX40 U51402 ( .A(\OFill[44][0] ), .B(n65641), .C(n65642), .D(n65643), .S0(
        n65814), .S1(N1082), .Q(n45588) );
  IMUX40 U51399 ( .A(\OFill[56][0] ), .B(n65621), .C(n65622), .D(n65623), .S0(
        n65802), .S1(n65923), .Q(n45581) );
  IMUX40 U51398 ( .A(\OFill[60][0] ), .B(n65625), .C(n65626), .D(n65627), .S0(
        n65784), .S1(n65538), .Q(n45583) );
  IMUX40 U51411 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65790), 
        .S1(n65922), .Q(n45596) );
  IMUX40 U51410 ( .A(n65672), .B(\OFill[13][0] ), .C(n65674), .D(n65675), .S0(
        n65809), .S1(n65922), .Q(n45598) );
  IMUX40 U62827 ( .A(n65636), .B(n65637), .C(\OFill[42][0] ), .D(n65639), .S0(
        n65823), .S1(n65921), .Q(n56466) );
  IMUX40 U62826 ( .A(n65640), .B(n65641), .C(\OFill[46][0] ), .D(n65643), .S0(
        n65822), .S1(n65914), .Q(n56468) );
  IMUX40 U62823 ( .A(n65620), .B(n65621), .C(\OFill[58][0] ), .D(n65623), .S0(
        n65828), .S1(N1256), .Q(n56461) );
  IMUX40 U62822 ( .A(n65624), .B(n65625), .C(\OFill[62][0] ), .D(n65627), .S0(
        n65820), .S1(N1112), .Q(n56463) );
  IMUX40 U62835 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(n65670), .D(n65671), 
        .S0(n65806), .S1(n65914), .Q(n56476) );
  IMUX40 U62834 ( .A(\OFill[12][0] ), .B(n65673), .C(\OFill[14][0] ), .D(
        n65675), .S0(n65804), .S1(n65914), .Q(n56478) );
  IMUX40 U62155 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65857), .S1(n65753), .Q(n55826) );
  IMUX40 U62154 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65873), .S1(n65752), .Q(n55828) );
  IMUX40 U62151 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65886), .S1(n65752), .Q(n55821) );
  IMUX40 U62150 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65887), .S1(n65752), .Q(n55823) );
  IMUX40 U62163 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65869), .S1(n65754), .Q(n55836) );
  IMUX40 U62162 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65869), .S1(n65755), .Q(n55838) );
  IMUX40 U63499 ( .A(n65636), .B(n65637), .C(\OFill[42][0] ), .D(n65639), .S0(
        n65895), .S1(n65778), .Q(n57106) );
  IMUX40 U63498 ( .A(n65640), .B(n65641), .C(\OFill[46][0] ), .D(n65643), .S0(
        n65899), .S1(n65760), .Q(n57108) );
  IMUX40 U63495 ( .A(n65620), .B(n65621), .C(\OFill[58][0] ), .D(n65623), .S0(
        n65888), .S1(n65759), .Q(n57101) );
  IMUX40 U63494 ( .A(n65624), .B(n65625), .C(\OFill[62][0] ), .D(n65627), .S0(
        n65879), .S1(n65759), .Q(n57103) );
  IMUX40 U63507 ( .A(n65668), .B(\OFill[9][0] ), .C(n65670), .D(n65671), .S0(
        n65863), .S1(n65772), .Q(n57116) );
  IMUX40 U63506 ( .A(n65672), .B(n65673), .C(\OFill[14][0] ), .D(n65675), .S0(
        n65859), .S1(n65776), .Q(n57118) );
  IMUX40 U64171 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65849), .S1(n65760), .Q(n57746) );
  IMUX40 U64170 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65908), .S1(n65762), .Q(n57748) );
  IMUX40 U64167 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65871), .S1(n65781), .Q(n57741) );
  IMUX40 U64166 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65896), .S1(n65780), .Q(n57743) );
  IMUX40 U64179 ( .A(n65668), .B(\OFill[9][0] ), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65865), .S1(n65759), .Q(n57756) );
  IMUX40 U64178 ( .A(n65672), .B(\OFill[13][0] ), .C(\OFill[14][0] ), .D(
        \OFill[15][0] ), .S0(n65901), .S1(n65774), .Q(n57758) );
  IMUX40 U65515 ( .A(n65636), .B(n65637), .C(\OFill[42][0] ), .D(
        \OFill[43][0] ), .S0(n65882), .S1(n65754), .Q(n59026) );
  IMUX40 U65514 ( .A(n65640), .B(n65641), .C(\OFill[46][0] ), .D(
        \OFill[47][0] ), .S0(n65891), .S1(n65749), .Q(n59028) );
  IMUX40 U65511 ( .A(n65620), .B(n65621), .C(\OFill[58][0] ), .D(
        \OFill[59][0] ), .S0(n65872), .S1(n65751), .Q(n59021) );
  IMUX40 U65510 ( .A(n65624), .B(n65625), .C(\OFill[62][0] ), .D(
        \OFill[63][0] ), .S0(n65860), .S1(n65750), .Q(n59023) );
  IMUX40 U65523 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65867), .S1(n65746), .Q(n59036) );
  IMUX40 U65522 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65878), .S1(n65753), .Q(n59038) );
  IMUX40 U17131 ( .A(\GFill[40][0] ), .B(n65701), .C(n65702), .D(n65703), .S0(
        n65897), .S1(n65747), .Q(n12946) );
  IMUX40 U17130 ( .A(\GFill[44][0] ), .B(n65705), .C(n65706), .D(n65707), .S0(
        n65902), .S1(n65748), .Q(n12948) );
  IMUX40 U17127 ( .A(\GFill[56][0] ), .B(n65685), .C(n65686), .D(n65687), .S0(
        n65900), .S1(n65744), .Q(n12941) );
  IMUX40 U17126 ( .A(\GFill[60][0] ), .B(n65689), .C(n65690), .D(n65691), .S0(
        n65902), .S1(n65746), .Q(n12943) );
  IMUX40 U17139 ( .A(\GFill[8][0] ), .B(n65733), .C(n65734), .D(n65735), .S0(
        n65883), .S1(n65750), .Q(n12956) );
  IMUX40 U17138 ( .A(\GFill[12][0] ), .B(n65737), .C(n65738), .D(n65739), .S0(
        n65858), .S1(n65752), .Q(n12958) );
  IMUX40 U16459 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65786), .S1(N1082), .Q(n12306) );
  IMUX40 U16458 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65786), .S1(n65923), .Q(n12308) );
  IMUX40 U16455 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65800), .S1(N1082), .Q(n12301) );
  IMUX40 U16454 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65819), .S1(n65538), .Q(n12303) );
  IMUX40 U16467 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65819), .S1(N1082), .Q(n12316) );
  IMUX40 U16466 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65816), .S1(n65538), .Q(n12318) );
  IMUX40 U18475 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65882), 
        .S1(n65781), .Q(n14226) );
  IMUX40 U18474 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65883), 
        .S1(n65776), .Q(n14228) );
  IMUX40 U18471 ( .A(\GFill[56][0] ), .B(n65685), .C(n65686), .D(n65687), .S0(
        n65847), .S1(n65769), .Q(n14221) );
  IMUX40 U18470 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(N1207), 
        .S1(n65765), .Q(n14223) );
  IMUX40 U18483 ( .A(n65732), .B(n65733), .C(n65734), .D(n65735), .S0(n65907), 
        .S1(n65780), .Q(n14236) );
  IMUX40 U18482 ( .A(n65736), .B(n65737), .C(n65738), .D(n65739), .S0(n65900), 
        .S1(n65781), .Q(n14238) );
  IMUX40 U17803 ( .A(n65700), .B(\GFill[41][0] ), .C(\GFill[42][0] ), .D(
        \GFill[43][0] ), .S0(n65837), .S1(n65745), .Q(n13586) );
  IMUX40 U17802 ( .A(n65704), .B(\GFill[45][0] ), .C(\GFill[46][0] ), .D(
        \GFill[47][0] ), .S0(n65837), .S1(n65755), .Q(n13588) );
  IMUX40 U17799 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65838), .S1(n65756), .Q(n13581) );
  IMUX40 U17798 ( .A(n65688), .B(\GFill[61][0] ), .C(\GFill[62][0] ), .D(
        \GFill[63][0] ), .S0(n65838), .S1(n65751), .Q(n13583) );
  IMUX40 U17811 ( .A(n65732), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(
        \GFill[11][0] ), .S0(n65834), .S1(N1208), .Q(n13596) );
  IMUX40 U17810 ( .A(n65736), .B(\GFill[13][0] ), .C(\GFill[14][0] ), .D(
        \GFill[15][0] ), .S0(n65834), .S1(n65745), .Q(n13598) );
  IMUX40 U19147 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(n65703), .S0(n65795), .S1(N1082), .Q(n14866) );
  IMUX40 U19146 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(n65707), .S0(n65819), .S1(n65923), .Q(n14868) );
  IMUX40 U19143 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(n65687), .S0(n65829), .S1(n65922), .Q(n14861) );
  IMUX40 U19142 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(n65691), .S0(n65786), .S1(N1082), .Q(n14863) );
  IMUX40 U19155 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(n65735), .S0(n65815), .S1(n65923), .Q(n14876) );
  IMUX40 U19154 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(n65739), .S0(n65822), .S1(n65922), .Q(n14878) );
  IMUX40 U30571 ( .A(n65700), .B(n65701), .C(\GFill[42][0] ), .D(n65703), .S0(
        n65830), .S1(n65921), .Q(n25746) );
  IMUX40 U30570 ( .A(n65704), .B(n65705), .C(\GFill[46][0] ), .D(n65707), .S0(
        n65821), .S1(n65914), .Q(n25748) );
  IMUX40 U30567 ( .A(n65684), .B(n65685), .C(\GFill[58][0] ), .D(n65687), .S0(
        n65830), .S1(N1184), .Q(n25741) );
  IMUX40 U30566 ( .A(n65688), .B(n65689), .C(\GFill[62][0] ), .D(n65691), .S0(
        n65831), .S1(N1172), .Q(n25743) );
  IMUX40 U30579 ( .A(n65732), .B(n65733), .C(\GFill[10][0] ), .D(n65735), .S0(
        n65789), .S1(n65913), .Q(n25756) );
  IMUX40 U30578 ( .A(n65736), .B(n65737), .C(\GFill[14][0] ), .D(n65739), .S0(
        n65782), .S1(N1112), .Q(n25758) );
  IMUX40 U29899 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65872), .S1(n65752), .Q(n25106) );
  IMUX40 U29898 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65877), .S1(n65752), .Q(n25108) );
  IMUX40 U29895 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65867), .S1(n65752), .Q(n25101) );
  IMUX40 U29894 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65833), .S1(n65752), .Q(n25103) );
  IMUX40 U29907 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65897), .S1(n65751), .Q(n25116) );
  IMUX40 U29906 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65908), .S1(n65750), .Q(n25118) );
  IMUX40 U31243 ( .A(n65700), .B(n65701), .C(\GFill[42][0] ), .D(n65703), .S0(
        n65870), .S1(n65759), .Q(n26386) );
  IMUX40 U31242 ( .A(n65704), .B(n65705), .C(\GFill[46][0] ), .D(n65707), .S0(
        n65853), .S1(n65781), .Q(n26388) );
  IMUX40 U31239 ( .A(n65684), .B(n65685), .C(\GFill[58][0] ), .D(n65687), .S0(
        N1207), .S1(n65759), .Q(n26381) );
  IMUX40 U31238 ( .A(n65688), .B(n65689), .C(\GFill[62][0] ), .D(n65691), .S0(
        n65858), .S1(n65759), .Q(n26383) );
  IMUX40 U31251 ( .A(n65732), .B(n65733), .C(\GFill[10][0] ), .D(n65735), .S0(
        n65894), .S1(n65775), .Q(n26396) );
  IMUX40 U31250 ( .A(n65736), .B(n65737), .C(\GFill[14][0] ), .D(n65739), .S0(
        n65893), .S1(n65760), .Q(n26398) );
  IMUX40 U32587 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65803), .S1(n65911), .Q(n27666) );
  IMUX40 U32586 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65785), .S1(n65922), .Q(n27668) );
  IMUX40 U32583 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65815), .S1(n65923), .Q(n27661) );
  IMUX40 U32582 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65827), .S1(N1082), .Q(n27663) );
  IMUX40 U32595 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65821), .S1(N1082), .Q(n27676) );
  IMUX40 U32594 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65801), .S1(N860), .Q(n27678) );
  IMUX40 U31915 ( .A(n65700), .B(n65701), .C(\GFill[42][0] ), .D(
        \GFill[43][0] ), .S0(n65910), .S1(n65766), .Q(n27026) );
  IMUX40 U31914 ( .A(n65704), .B(n65705), .C(\GFill[46][0] ), .D(
        \GFill[47][0] ), .S0(n65893), .S1(n65762), .Q(n27028) );
  IMUX40 U31911 ( .A(n65684), .B(n65685), .C(\GFill[58][0] ), .D(
        \GFill[59][0] ), .S0(n65898), .S1(n65764), .Q(n27021) );
  IMUX40 U31910 ( .A(n65688), .B(n65689), .C(\GFill[62][0] ), .D(
        \GFill[63][0] ), .S0(n65841), .S1(n65760), .Q(n27023) );
  IMUX40 U31923 ( .A(n65732), .B(n65733), .C(\GFill[10][0] ), .D(
        \GFill[11][0] ), .S0(n65837), .S1(n65767), .Q(n27036) );
  IMUX40 U31922 ( .A(n65736), .B(n65737), .C(\GFill[14][0] ), .D(
        \GFill[15][0] ), .S0(n65881), .S1(n65766), .Q(n27038) );
  IMUX40 U33259 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(n65703), .S0(n65864), .S1(n65744), .Q(n28306) );
  IMUX40 U33258 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(n65707), .S0(n65833), .S1(N1208), .Q(n28308) );
  IMUX40 U33255 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(n65687), .S0(n65876), .S1(n65746), .Q(n28301) );
  IMUX40 U33254 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(n65691), .S0(n65902), .S1(n65757), .Q(n28303) );
  IMUX40 U33267 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(n65735), .S0(n65889), .S1(n65744), .Q(n28316) );
  IMUX40 U33266 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(n65739), .S0(n65875), .S1(n65744), .Q(n28318) );
  IMUX40 U23179 ( .A(n65700), .B(n65701), .C(n65702), .D(\GFill[43][0] ), .S0(
        n65843), .S1(n65754), .Q(n18706) );
  IMUX40 U23178 ( .A(n65704), .B(n65705), .C(n65706), .D(\GFill[47][0] ), .S0(
        n65881), .S1(n65753), .Q(n18708) );
  IMUX40 U23175 ( .A(\GFill[56][0] ), .B(n65685), .C(n65686), .D(
        \GFill[59][0] ), .S0(n65852), .S1(n65752), .Q(n18701) );
  IMUX40 U23174 ( .A(n65688), .B(n65689), .C(n65690), .D(\GFill[63][0] ), .S0(
        n65867), .S1(n65753), .Q(n18703) );
  IMUX40 U23187 ( .A(n65732), .B(n65733), .C(n65734), .D(\GFill[11][0] ), .S0(
        n65878), .S1(n65752), .Q(n18716) );
  IMUX40 U23186 ( .A(n65736), .B(n65737), .C(n65738), .D(\GFill[15][0] ), .S0(
        n65839), .S1(N1208), .Q(n18718) );
  IMUX40 U22507 ( .A(\GFill[40][0] ), .B(n65701), .C(n65702), .D(
        \GFill[43][0] ), .S0(n65796), .S1(n65914), .Q(n18066) );
  IMUX40 U22506 ( .A(\GFill[44][0] ), .B(n65705), .C(n65706), .D(
        \GFill[47][0] ), .S0(n65794), .S1(n65921), .Q(n18068) );
  IMUX40 U22503 ( .A(\GFill[56][0] ), .B(n65685), .C(n65686), .D(
        \GFill[59][0] ), .S0(n65805), .S1(n65914), .Q(n18061) );
  IMUX40 U22502 ( .A(\GFill[60][0] ), .B(n65689), .C(n65690), .D(
        \GFill[63][0] ), .S0(n65800), .S1(n65921), .Q(n18063) );
  IMUX40 U22515 ( .A(\GFill[8][0] ), .B(n65733), .C(n65734), .D(\GFill[11][0] ), .S0(n65828), .S1(n65914), .Q(n18076) );
  IMUX40 U22514 ( .A(\GFill[12][0] ), .B(n65737), .C(n65738), .D(
        \GFill[15][0] ), .S0(n65807), .S1(n65913), .Q(n18078) );
  IMUX40 U35275 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65834), 
        .S1(n65754), .Q(n30226) );
  IMUX40 U35274 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65880), 
        .S1(n65754), .Q(n30228) );
  IMUX40 U35271 ( .A(n65684), .B(n65685), .C(n65686), .D(n65687), .S0(n65905), 
        .S1(n65754), .Q(n30221) );
  IMUX40 U35270 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(n65881), 
        .S1(n65754), .Q(n30223) );
  IMUX40 U54091 ( .A(n65636), .B(\OFill[41][0] ), .C(\OFill[42][0] ), .D(
        \OFill[43][0] ), .S0(n65851), .S1(n65774), .Q(n48146) );
  IMUX40 U54090 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65851), .S1(n65774), .Q(n48148) );
  IMUX40 U54087 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65850), .S1(n65780), .Q(n48141) );
  IMUX40 U54086 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65850), .S1(n65763), .Q(n48143) );
  IMUX40 U54099 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65865), .S1(n65764), .Q(n48156) );
  IMUX40 U54098 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65863), .S1(n65781), .Q(n48158) );
  IMUX40 U55435 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(n65639), .S0(n65890), .S1(n65749), .Q(n49426) );
  IMUX40 U55434 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(n65643), .S0(n65840), .S1(N1208), .Q(n49428) );
  IMUX40 U55431 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(n65623), .S0(n65856), .S1(n65755), .Q(n49421) );
  IMUX40 U55430 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(n65627), .S0(n65858), .S1(N1208), .Q(n49423) );
  IMUX40 U55443 ( .A(n65668), .B(\OFill[9][0] ), .C(n65670), .D(n65671), .S0(
        n65866), .S1(n65749), .Q(n49436) );
  IMUX40 U55442 ( .A(n65672), .B(\OFill[13][0] ), .C(n65674), .D(n65675), .S0(
        n65867), .S1(n65749), .Q(n49438) );
  IMUX40 U67531 ( .A(\OFill[40][0] ), .B(n65637), .C(n65638), .D(n65639), .S0(
        n65850), .S1(n65747), .Q(n60946) );
  IMUX40 U67530 ( .A(\OFill[44][0] ), .B(n65641), .C(n65642), .D(n65643), .S0(
        N1207), .S1(n65747), .Q(n60948) );
  IMUX40 U67527 ( .A(\OFill[56][0] ), .B(n65621), .C(n65622), .D(n65623), .S0(
        n65892), .S1(n65747), .Q(n60941) );
  IMUX40 U67526 ( .A(\OFill[60][0] ), .B(n65625), .C(n65626), .D(n65627), .S0(
        n65902), .S1(n65747), .Q(n60943) );
  IMUX40 U9067 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(n65702), .D(
        \GFill[43][0] ), .S0(n65789), .S1(N704), .Q(n5266) );
  IMUX40 U9066 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(n65706), .D(
        \GFill[47][0] ), .S0(n65782), .S1(N704), .Q(n5268) );
  IMUX40 U9063 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(n65686), .D(
        \GFill[59][0] ), .S0(n65809), .S1(N704), .Q(n5261) );
  IMUX40 U9062 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(n65690), .D(
        \GFill[63][0] ), .S0(n65817), .S1(N704), .Q(n5263) );
  IMUX40 U8395 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65809), .S1(n65536), .Q(n4626) );
  IMUX40 U8394 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65809), .S1(n65536), .Q(n4628) );
  IMUX40 U8391 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65810), .S1(n65536), .Q(n4621) );
  IMUX40 U8390 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65810), .S1(n65536), .Q(n4623) );
  IMUX40 U8403 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(n65734), .D(
        \GFill[11][0] ), .S0(n65789), .S1(n65536), .Q(n4636) );
  IMUX40 U8402 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(n65738), .D(
        \GFill[15][0] ), .S0(n65789), .S1(n65536), .Q(n4638) );
  IMUX40 U10411 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(n65702), .D(
        \GFill[43][0] ), .S0(n65819), .S1(N716), .Q(n6546) );
  IMUX40 U10410 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(n65706), .D(
        \GFill[47][0] ), .S0(n65819), .S1(N716), .Q(n6548) );
  IMUX40 U10407 ( .A(n65684), .B(\GFill[57][0] ), .C(n65686), .D(
        \GFill[59][0] ), .S0(n65819), .S1(N716), .Q(n6541) );
  IMUX40 U10406 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(n65690), .D(
        \GFill[63][0] ), .S0(n65819), .S1(N716), .Q(n6543) );
  IMUX40 U9739 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65800), .S1(n65935), .Q(n5906) );
  IMUX40 U9738 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65799), .S1(n65934), .Q(n5908) );
  IMUX40 U9735 ( .A(n65684), .B(\GFill[57][0] ), .C(\GFill[58][0] ), .D(
        \GFill[59][0] ), .S0(n65799), .S1(n65934), .Q(n5901) );
  IMUX40 U9734 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65799), .S1(n65935), .Q(n5903) );
  IMUX40 U9747 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(
        \GFill[11][0] ), .S0(n65798), .S1(n65935), .Q(n5916) );
  IMUX40 U9746 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65798), .S1(n65935), .Q(n5918) );
  IMUX40 U11083 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(n65702), .D(
        \GFill[43][0] ), .S0(n65830), .S1(N722), .Q(n7186) );
  IMUX40 U11082 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(n65706), .D(
        \GFill[47][0] ), .S0(n65830), .S1(N722), .Q(n7188) );
  IMUX40 U11079 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(n65686), .D(
        \GFill[59][0] ), .S0(n65830), .S1(N722), .Q(n7181) );
  IMUX40 U11078 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(n65690), .D(
        \GFill[63][0] ), .S0(n65829), .S1(N722), .Q(n7183) );
  IMUX40 U12427 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65804), .S1(n65933), .Q(n8466) );
  IMUX40 U12426 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65804), .S1(N1022), .Q(n8468) );
  IMUX40 U12423 ( .A(n65684), .B(\GFill[57][0] ), .C(\GFill[58][0] ), .D(
        \GFill[59][0] ), .S0(n65804), .S1(n65930), .Q(n8461) );
  IMUX40 U12422 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65804), .S1(n65932), .Q(n8463) );
  IMUX40 U12435 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(n65734), .D(
        \GFill[11][0] ), .S0(n65803), .S1(n65930), .Q(n8476) );
  IMUX40 U12434 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(n65738), .D(
        \GFill[15][0] ), .S0(n65802), .S1(n65932), .Q(n8478) );
  IMUX40 U13771 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65791), .S1(n65929), .Q(n9746) );
  IMUX40 U13770 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65791), .S1(n65928), .Q(n9748) );
  IMUX40 U13767 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65791), .S1(n65928), .Q(n9741) );
  IMUX40 U13766 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65791), .S1(n65929), .Q(n9743) );
  IMUX40 U13779 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65790), .S1(n65929), .Q(n9756) );
  IMUX40 U13778 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65790), .S1(n65929), .Q(n9758) );
  IMUX40 U15115 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65796), .S1(N1010), .Q(n11026) );
  IMUX40 U15114 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65796), .S1(n65925), .Q(n11028) );
  IMUX40 U15111 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65795), .S1(n65925), .Q(n11021) );
  IMUX40 U15110 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65795), .S1(n65924), .Q(n11023) );
  IMUX40 U15123 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(n65734), .D(
        \GFill[11][0] ), .S0(n65794), .S1(N1010), .Q(n11036) );
  IMUX40 U15122 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(n65738), .D(
        \GFill[15][0] ), .S0(n65794), .S1(n65925), .Q(n11038) );
  IMUX40 U14443 ( .A(n65700), .B(\GFill[41][0] ), .C(\GFill[42][0] ), .D(
        n65703), .S0(n65807), .S1(n65927), .Q(n10386) );
  IMUX40 U14442 ( .A(n65704), .B(\GFill[45][0] ), .C(\GFill[46][0] ), .D(
        n65707), .S0(n65807), .S1(n65926), .Q(n10388) );
  IMUX40 U14439 ( .A(n65684), .B(\GFill[57][0] ), .C(\GFill[58][0] ), .D(
        n65687), .S0(n65807), .S1(n65926), .Q(n10381) );
  IMUX40 U14438 ( .A(n65688), .B(\GFill[61][0] ), .C(\GFill[62][0] ), .D(
        n65691), .S0(n65807), .S1(n65927), .Q(n10383) );
  IMUX40 U14451 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65802), .S1(n65927), .Q(n10396) );
  IMUX40 U14450 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65798), .S1(n65927), .Q(n10398) );
  IMUX40 U27883 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(n65703), .S0(n65906), .S1(n65772), .Q(n23186) );
  IMUX40 U27882 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(n65707), .S0(n65907), .S1(n65772), .Q(n23188) );
  IMUX40 U27879 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(n65687), .S0(n65888), .S1(n65777), .Q(n23181) );
  IMUX40 U27878 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(n65691), .S0(n65889), .S1(n65771), .Q(n23183) );
  IMUX40 U29227 ( .A(n65700), .B(\GFill[41][0] ), .C(\GFill[42][0] ), .D(
        \GFill[43][0] ), .S0(n65795), .S1(n65921), .Q(n24466) );
  IMUX40 U29226 ( .A(n65704), .B(\GFill[45][0] ), .C(\GFill[46][0] ), .D(
        \GFill[47][0] ), .S0(n65797), .S1(n65914), .Q(n24468) );
  IMUX40 U29223 ( .A(n65684), .B(\GFill[57][0] ), .C(\GFill[58][0] ), .D(
        \GFill[59][0] ), .S0(n65790), .S1(n65921), .Q(n24461) );
  IMUX40 U29222 ( .A(n65688), .B(\GFill[61][0] ), .C(\GFill[62][0] ), .D(
        \GFill[63][0] ), .S0(n65831), .S1(n65914), .Q(n24463) );
  IMUX40 U29235 ( .A(n65732), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(n65735), .S0(n65803), .S1(N1184), .Q(n24476) );
  IMUX40 U29234 ( .A(n65736), .B(\GFill[13][0] ), .C(\GFill[14][0] ), .D(
        n65739), .S0(n65821), .S1(n65921), .Q(n24478) );
  IMUX40 U25867 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(n65703), .S0(n65892), .S1(n65778), .Q(n21266) );
  IMUX40 U25866 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(n65707), .S0(n65888), .S1(n65779), .Q(n21268) );
  IMUX40 U25863 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(n65687), .S0(n65845), .S1(n65781), .Q(n21261) );
  IMUX40 U25862 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(n65691), .S0(n65837), .S1(n65779), .Q(n21263) );
  IMUX40 U27211 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65905), .S1(n65746), .Q(n22546) );
  IMUX40 U27210 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65842), .S1(n65745), .Q(n22548) );
  IMUX40 U27207 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65864), .S1(n65745), .Q(n22541) );
  IMUX40 U27206 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65847), .S1(n65745), .Q(n22543) );
  IMUX40 U27219 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65896), .S1(n65746), .Q(n22556) );
  IMUX40 U27218 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65873), .S1(n65746), .Q(n22558) );
  IMUX40 U24523 ( .A(n65700), .B(\GFill[41][0] ), .C(\GFill[42][0] ), .D(
        \GFill[43][0] ), .S0(n65805), .S1(N842), .Q(n19986) );
  IMUX40 U24522 ( .A(n65704), .B(\GFill[45][0] ), .C(\GFill[46][0] ), .D(
        \GFill[47][0] ), .S0(n65831), .S1(N842), .Q(n19988) );
  IMUX40 U24519 ( .A(n65684), .B(\GFill[57][0] ), .C(\GFill[58][0] ), .D(
        \GFill[59][0] ), .S0(n65786), .S1(N842), .Q(n19981) );
  IMUX40 U24518 ( .A(n65688), .B(\GFill[61][0] ), .C(\GFill[62][0] ), .D(
        \GFill[63][0] ), .S0(n65830), .S1(N842), .Q(n19983) );
  IMUX40 U24531 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65817), .S1(N842), .Q(n19996) );
  IMUX40 U24530 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65786), .S1(N842), .Q(n19998) );
  IMUX40 U23851 ( .A(\GFill[40][0] ), .B(n65701), .C(n65702), .D(
        \GFill[43][0] ), .S0(n65839), .S1(n65780), .Q(n19346) );
  IMUX40 U23850 ( .A(\GFill[44][0] ), .B(n65705), .C(n65706), .D(
        \GFill[47][0] ), .S0(n65871), .S1(n65775), .Q(n19348) );
  IMUX40 U23847 ( .A(\GFill[56][0] ), .B(n65685), .C(n65686), .D(
        \GFill[59][0] ), .S0(n65849), .S1(n65767), .Q(n19341) );
  IMUX40 U23846 ( .A(\GFill[60][0] ), .B(n65689), .C(n65690), .D(
        \GFill[63][0] ), .S0(n65852), .S1(n65765), .Q(n19343) );
  IMUX40 U23859 ( .A(n65732), .B(n65733), .C(n65734), .D(\GFill[11][0] ), .S0(
        n65889), .S1(n65765), .Q(n19356) );
  IMUX40 U23858 ( .A(n65736), .B(n65737), .C(n65738), .D(\GFill[15][0] ), .S0(
        N1207), .S1(n65779), .Q(n19358) );
  IMUX40 U41323 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(n65638), .D(
        \OFill[43][0] ), .S0(n65816), .S1(n65929), .Q(n35986) );
  IMUX40 U41322 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(n65642), .D(
        \OFill[47][0] ), .S0(n65817), .S1(N1004), .Q(n35988) );
  IMUX40 U41319 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(n65622), .D(
        \OFill[59][0] ), .S0(n65817), .S1(N1004), .Q(n35981) );
  IMUX40 U41318 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(n65626), .D(
        \OFill[63][0] ), .S0(n65817), .S1(N1004), .Q(n35983) );
  IMUX40 U42667 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65828), .S1(N1034), .Q(n37266) );
  IMUX40 U42666 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65828), .S1(N1034), .Q(n37268) );
  IMUX40 U42663 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65827), .S1(N1034), .Q(n37261) );
  IMUX40 U42662 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65827), .S1(N1034), .Q(n37263) );
  IMUX40 U41995 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(n65638), .D(
        \OFill[43][0] ), .S0(n65802), .S1(n65934), .Q(n36626) );
  IMUX40 U41994 ( .A(n65640), .B(\OFill[45][0] ), .C(n65642), .D(
        \OFill[47][0] ), .S0(n65802), .S1(n65935), .Q(n36628) );
  IMUX40 U41991 ( .A(n65620), .B(\OFill[57][0] ), .C(n65622), .D(
        \OFill[59][0] ), .S0(n65799), .S1(n65934), .Q(n36621) );
  IMUX40 U41990 ( .A(n65624), .B(\OFill[61][0] ), .C(n65626), .D(
        \OFill[63][0] ), .S0(n65799), .S1(n65935), .Q(n36623) );
  IMUX40 U42003 ( .A(\OFill[8][0] ), .B(n65669), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65800), .S1(n65934), .Q(n36636) );
  IMUX40 U42002 ( .A(\OFill[12][0] ), .B(n65673), .C(n65674), .D(
        \OFill[15][0] ), .S0(n65800), .S1(n65934), .Q(n36638) );
  IMUX40 U43339 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65826), .S1(N1010), .Q(n37906) );
  IMUX40 U43338 ( .A(n65640), .B(\OFill[45][0] ), .C(\OFill[46][0] ), .D(
        \OFill[47][0] ), .S0(n65825), .S1(N980), .Q(n37908) );
  IMUX40 U43335 ( .A(n65620), .B(\OFill[57][0] ), .C(\OFill[58][0] ), .D(
        \OFill[59][0] ), .S0(n65825), .S1(n65925), .Q(n37901) );
  IMUX40 U43334 ( .A(n65624), .B(\OFill[61][0] ), .C(\OFill[62][0] ), .D(
        \OFill[63][0] ), .S0(n65825), .S1(n65924), .Q(n37903) );
  IMUX40 U44683 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(n65638), .D(
        \OFill[43][0] ), .S0(n65806), .S1(n65933), .Q(n39186) );
  IMUX40 U44682 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(n65642), .D(
        \OFill[47][0] ), .S0(n65806), .S1(n65930), .Q(n39188) );
  IMUX40 U44679 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(n65622), .D(
        \OFill[59][0] ), .S0(n65803), .S1(n65932), .Q(n39181) );
  IMUX40 U44678 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(n65626), .D(
        \OFill[63][0] ), .S0(n65803), .S1(n65933), .Q(n39183) );
  IMUX40 U44691 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65805), .S1(n65931), .Q(n39196) );
  IMUX40 U44690 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65805), .S1(n65933), .Q(n39198) );
  IMUX40 U45355 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65821), .S1(N1040), .Q(n39826) );
  IMUX40 U45354 ( .A(n65640), .B(\OFill[45][0] ), .C(\OFill[46][0] ), .D(
        \OFill[47][0] ), .S0(n65821), .S1(N1040), .Q(n39828) );
  IMUX40 U45351 ( .A(n65620), .B(\OFill[57][0] ), .C(\OFill[58][0] ), .D(
        \OFill[59][0] ), .S0(n65820), .S1(N1040), .Q(n39821) );
  IMUX40 U45350 ( .A(n65624), .B(\OFill[61][0] ), .C(\OFill[62][0] ), .D(
        \OFill[63][0] ), .S0(n65820), .S1(N1040), .Q(n39823) );
  IMUX40 U46695 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65799), .S1(n65926), .Q(n41101) );
  IMUX40 U46694 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65807), .S1(n65927), .Q(n41103) );
  IMUX40 U46707 ( .A(\OFill[8][0] ), .B(n65669), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65807), .S1(n65926), .Q(n41116) );
  IMUX40 U46706 ( .A(\OFill[12][0] ), .B(n65673), .C(n65674), .D(
        \OFill[15][0] ), .S0(n65818), .S1(n65926), .Q(n41118) );
  IMUX40 U46027 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65793), .S1(n65928), .Q(n40466) );
  IMUX40 U46026 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65793), .S1(n65929), .Q(n40468) );
  IMUX40 U46023 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65790), .S1(n65928), .Q(n40461) );
  IMUX40 U46022 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65791), .S1(n65929), .Q(n40463) );
  IMUX40 U46035 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65792), .S1(n65928), .Q(n40476) );
  IMUX40 U46034 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65792), .S1(n65928), .Q(n40478) );
  IMUX40 U47371 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65814), .S1(N1010), .Q(n41746) );
  IMUX40 U47370 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65815), .S1(n65925), .Q(n41748) );
  IMUX40 U47367 ( .A(n65620), .B(\OFill[57][0] ), .C(\OFill[58][0] ), .D(
        n65623), .S0(n65795), .S1(n65924), .Q(n41741) );
  IMUX40 U47366 ( .A(n65624), .B(\OFill[61][0] ), .C(\OFill[62][0] ), .D(
        n65627), .S0(n65795), .S1(N1010), .Q(n41743) );
  IMUX40 U47379 ( .A(\OFill[8][0] ), .B(n65669), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65797), .S1(n65924), .Q(n41756) );
  IMUX40 U47378 ( .A(\OFill[12][0] ), .B(n65673), .C(\OFill[14][0] ), .D(
        \OFill[15][0] ), .S0(n65797), .S1(n65924), .Q(n41758) );
  IMUX40 U60139 ( .A(n65636), .B(\OFill[41][0] ), .C(\OFill[42][0] ), .D(
        n65639), .S0(n65867), .S1(n65770), .Q(n53906) );
  IMUX40 U60138 ( .A(n65640), .B(\OFill[45][0] ), .C(\OFill[46][0] ), .D(
        n65643), .S0(n65853), .S1(n65770), .Q(n53908) );
  IMUX40 U60135 ( .A(n65620), .B(\OFill[57][0] ), .C(\OFill[58][0] ), .D(
        n65623), .S0(n65879), .S1(n65770), .Q(n53901) );
  IMUX40 U60134 ( .A(n65624), .B(\OFill[61][0] ), .C(\OFill[62][0] ), .D(
        n65627), .S0(n65903), .S1(n65770), .Q(n53903) );
  IMUX40 U61483 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(n65639), .S0(n65828), .S1(n65914), .Q(n55186) );
  IMUX40 U61482 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(n65643), .S0(n65820), .S1(n65913), .Q(n55188) );
  IMUX40 U61479 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(n65623), .S0(n65830), .S1(n65914), .Q(n55181) );
  IMUX40 U61478 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(n65627), .S0(n65789), .S1(N1172), .Q(n55183) );
  IMUX40 U61491 ( .A(n65668), .B(\OFill[9][0] ), .C(n65670), .D(n65671), .S0(
        n65800), .S1(n65914), .Q(n55196) );
  IMUX40 U61490 ( .A(n65672), .B(n65673), .C(\OFill[14][0] ), .D(n65675), .S0(
        n65786), .S1(N1112), .Q(n55198) );
  IMUX40 U58123 ( .A(n65636), .B(\OFill[41][0] ), .C(\OFill[42][0] ), .D(
        \OFill[43][0] ), .S0(n65898), .S1(n65773), .Q(n51986) );
  IMUX40 U58122 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65880), .S1(n65768), .Q(n51988) );
  IMUX40 U58119 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65905), .S1(n65767), .Q(n51981) );
  IMUX40 U58118 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65863), .S1(n65766), .Q(n51983) );
  IMUX40 U59467 ( .A(n65636), .B(\OFill[41][0] ), .C(\OFill[42][0] ), .D(
        n65639), .S0(n65883), .S1(n65745), .Q(n53266) );
  IMUX40 U59466 ( .A(n65640), .B(\OFill[45][0] ), .C(\OFill[46][0] ), .D(
        n65643), .S0(n65882), .S1(n65745), .Q(n53268) );
  IMUX40 U59463 ( .A(n65620), .B(\OFill[57][0] ), .C(\OFill[58][0] ), .D(
        n65623), .S0(n65851), .S1(n65745), .Q(n53261) );
  IMUX40 U59462 ( .A(n65624), .B(\OFill[61][0] ), .C(\OFill[62][0] ), .D(
        n65627), .S0(n65850), .S1(n65745), .Q(n53263) );
  IMUX40 U59475 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(n65670), .D(n65671), 
        .S0(n65882), .S1(n65744), .Q(n53276) );
  IMUX40 U59474 ( .A(\OFill[12][0] ), .B(n65673), .C(\OFill[14][0] ), .D(
        n65675), .S0(n65875), .S1(n65744), .Q(n53278) );
  IMUX40 U56107 ( .A(\OFill[40][0] ), .B(n65637), .C(n65638), .D(
        \OFill[43][0] ), .S0(n65855), .S1(n65774), .Q(n50066) );
  IMUX40 U56106 ( .A(\OFill[44][0] ), .B(n65641), .C(n65642), .D(
        \OFill[47][0] ), .S0(n65886), .S1(n65774), .Q(n50068) );
  IMUX40 U56103 ( .A(\OFill[56][0] ), .B(n65621), .C(n65622), .D(
        \OFill[59][0] ), .S0(n65849), .S1(n65777), .Q(n50061) );
  IMUX40 U56102 ( .A(\OFill[60][0] ), .B(n65625), .C(n65626), .D(
        \OFill[63][0] ), .S0(n65833), .S1(n65779), .Q(n50063) );
  IMUX40 U57451 ( .A(\OFill[40][0] ), .B(n65637), .C(n65638), .D(
        \OFill[43][0] ), .S0(n65904), .S1(n65748), .Q(n51346) );
  IMUX40 U57450 ( .A(\OFill[44][0] ), .B(n65641), .C(n65642), .D(
        \OFill[47][0] ), .S0(n65899), .S1(n65748), .Q(n51348) );
  IMUX40 U57447 ( .A(\OFill[56][0] ), .B(n65621), .C(n65622), .D(
        \OFill[59][0] ), .S0(n65886), .S1(n65749), .Q(n51341) );
  IMUX40 U57446 ( .A(\OFill[60][0] ), .B(n65625), .C(n65626), .D(
        \OFill[63][0] ), .S0(n65858), .S1(n65749), .Q(n51343) );
  IMUX40 U37291 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65827), 
        .S1(N956), .Q(n32146) );
  IMUX40 U37290 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65819), 
        .S1(N956), .Q(n32148) );
  IMUX40 U37287 ( .A(n65684), .B(n65685), .C(n65686), .D(n65687), .S0(n65805), 
        .S1(N956), .Q(n32141) );
  IMUX40 U37286 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(n65795), 
        .S1(N956), .Q(n32143) );
  IMUX40 U37295 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65790), 
        .S1(N956), .Q(n32151) );
  IMUX40 U37294 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65795), 
        .S1(N956), .Q(n32153) );
  IMUX40 U44018 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(n65674), .D(
        \OFill[15][0] ), .S0(n65819), .S1(n65931), .Q(n38558) );
  IMUX40 U69551 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65791), 
        .S1(N1244), .Q(n62871) );
  IMUX40 U69550 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65784), 
        .S1(N1244), .Q(n62873) );
  IMUX40 U11755 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65812), .S1(n65931), .Q(n7826) );
  IMUX40 U11754 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65810), .S1(n65931), .Q(n7828) );
  IMUX40 U11751 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65812), .S1(n65932), .Q(n7821) );
  IMUX40 U11750 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65790), .S1(n65931), .Q(n7823) );
  IMUX40 U11763 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65791), .S1(n65933), .Q(n7836) );
  IMUX40 U11762 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65790), .S1(n65930), .Q(n7838) );
  IMUX40 U38635 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65818), 
        .S1(N968), .Q(n33426) );
  IMUX40 U38634 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65784), 
        .S1(N968), .Q(n33428) );
  IMUX40 U38631 ( .A(n65684), .B(n65685), .C(n65686), .D(n65687), .S0(n65810), 
        .S1(N968), .Q(n33421) );
  IMUX40 U38630 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(n65810), 
        .S1(N968), .Q(n33423) );
  IMUX40 U38643 ( .A(n65732), .B(n65733), .C(n65734), .D(n65735), .S0(n65826), 
        .S1(N968), .Q(n33436) );
  IMUX40 U38642 ( .A(n65736), .B(n65737), .C(n65738), .D(n65739), .S0(n65825), 
        .S1(N968), .Q(n33438) );
  IMUX40 U44011 ( .A(n65636), .B(\OFill[41][0] ), .C(\OFill[42][0] ), .D(
        n65639), .S0(n65824), .S1(n65933), .Q(n38546) );
  IMUX40 U44010 ( .A(n65640), .B(\OFill[45][0] ), .C(\OFill[46][0] ), .D(
        n65643), .S0(n65823), .S1(n65930), .Q(n38548) );
  IMUX40 U44007 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65818), .S1(n65930), .Q(n38541) );
  IMUX40 U44006 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65827), .S1(n65932), .Q(n38543) );
  IMUX40 U44019 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65811), .S1(n65931), .Q(n38556) );
  IMUX40 U46699 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65782), .S1(n65926), .Q(n41106) );
  IMUX40 U46698 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65782), .S1(n65927), .Q(n41108) );
  IMUX40 U69547 ( .A(n65636), .B(n65637), .C(n65638), .D(n65639), .S0(n65803), 
        .S1(N1244), .Q(n62866) );
  IMUX40 U69546 ( .A(n65640), .B(n65641), .C(n65642), .D(n65643), .S0(n65797), 
        .S1(N1244), .Q(n62868) );
  IMUX40 U69543 ( .A(n65620), .B(n65621), .C(n65622), .D(n65623), .S0(n65806), 
        .S1(N1244), .Q(n62861) );
  IMUX40 U69542 ( .A(n65624), .B(n65625), .C(n65626), .D(n65627), .S0(n65829), 
        .S1(N1244), .Q(n62863) );
  IMUX40 U25197 ( .A(\GFill[32][0] ), .B(n65693), .C(n65694), .D(n65695), .S0(
        n65893), .S1(n65749), .Q(n20625) );
  IMUX40 U25194 ( .A(n65704), .B(\GFill[45][0] ), .C(\GFill[46][0] ), .D(
        \GFill[47][0] ), .S0(n65855), .S1(n65752), .Q(n20628) );
  IMUX40 U25195 ( .A(n65700), .B(\GFill[41][0] ), .C(\GFill[42][0] ), .D(
        \GFill[43][0] ), .S0(n65910), .S1(n65754), .Q(n20626) );
  IMUX40 U25031 ( .A(n20625), .B(n20626), .C(n20627), .D(n20628), .S0(N850), 
        .S1(n65920), .Q(n20624) );
  IMUX40 U25193 ( .A(\GFill[48][0] ), .B(n65677), .C(n65678), .D(n65679), .S0(
        n65855), .S1(n65751), .Q(n20620) );
  IMUX40 U25190 ( .A(n65688), .B(\GFill[61][0] ), .C(\GFill[62][0] ), .D(
        \GFill[63][0] ), .S0(n65854), .S1(n65756), .Q(n20623) );
  IMUX40 U25191 ( .A(n65684), .B(\GFill[57][0] ), .C(\GFill[58][0] ), .D(
        \GFill[59][0] ), .S0(n65854), .S1(n65754), .Q(n20621) );
  IMUX40 U25030 ( .A(n20620), .B(n20621), .C(n20622), .D(n20623), .S0(N850), 
        .S1(n65920), .Q(n20619) );
  IMUX40 U54765 ( .A(\OFill[32][0] ), .B(n65629), .C(n65630), .D(n65631), .S0(
        n65810), .S1(n65913), .Q(n48785) );
  IMUX40 U54762 ( .A(n65640), .B(\OFill[45][0] ), .C(\OFill[46][0] ), .D(
        \OFill[47][0] ), .S0(n65782), .S1(N1112), .Q(n48788) );
  IMUX40 U54763 ( .A(n65636), .B(\OFill[41][0] ), .C(\OFill[42][0] ), .D(
        \OFill[43][0] ), .S0(n65789), .S1(n65913), .Q(n48786) );
  IMUX40 U54599 ( .A(n48785), .B(n48786), .C(n48787), .D(n48788), .S0(N1114), 
        .S1(N1113), .Q(n48784) );
  IMUX40 U54761 ( .A(\OFill[48][0] ), .B(n65613), .C(n65614), .D(n65615), .S0(
        n65787), .S1(N1112), .Q(n48780) );
  IMUX40 U54758 ( .A(n65624), .B(\OFill[61][0] ), .C(\OFill[62][0] ), .D(
        \OFill[63][0] ), .S0(n65808), .S1(N1184), .Q(n48783) );
  IMUX40 U54759 ( .A(n65620), .B(\OFill[57][0] ), .C(\OFill[58][0] ), .D(
        \OFill[59][0] ), .S0(n65817), .S1(n65913), .Q(n48781) );
  IMUX40 U54598 ( .A(n48780), .B(n48781), .C(n48782), .D(n48783), .S0(N1114), 
        .S1(N1113), .Q(n48779) );
  IMUX40 U7725 ( .A(\GFill[32][0] ), .B(n65693), .C(\GFill[34][0] ), .D(n65695), .S0(n65787), .S1(n65535), .Q(n3985) );
  IMUX40 U7722 ( .A(n65704), .B(n65705), .C(\GFill[46][0] ), .D(n65707), .S0(
        n65788), .S1(n65535), .Q(n3988) );
  IMUX40 U7723 ( .A(n65700), .B(n65701), .C(\GFill[42][0] ), .D(n65703), .S0(
        n65788), .S1(n65535), .Q(n3986) );
  IMUX40 U7559 ( .A(n3985), .B(n3986), .C(n3987), .D(n3988), .S0(N694), .S1(
        N693), .Q(n3984) );
  IMUX40 U7721 ( .A(\GFill[48][0] ), .B(n65677), .C(\GFill[50][0] ), .D(n65679), .S0(n65788), .S1(n65535), .Q(n3980) );
  IMUX40 U7718 ( .A(n65688), .B(n65689), .C(\GFill[62][0] ), .D(n65691), .S0(
        n65788), .S1(n65535), .Q(n3983) );
  IMUX40 U7719 ( .A(n65684), .B(n65685), .C(\GFill[58][0] ), .D(n65687), .S0(
        n65788), .S1(n65535), .Q(n3981) );
  IMUX40 U7558 ( .A(n3980), .B(n3981), .C(n3982), .D(n3983), .S0(N694), .S1(
        N693), .Q(n3979) );
  IMUX40 U37965 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(n65876), 
        .S1(N1208), .Q(n32785) );
  IMUX40 U37961 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65878), 
        .S1(n65746), .Q(n32780) );
  IMUX40 U35949 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(n65863), 
        .S1(n65764), .Q(n30865) );
  IMUX40 U35945 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65874), 
        .S1(n65765), .Q(n30860) );
  IMUX40 U35957 ( .A(n65724), .B(n65725), .C(n65726), .D(n65727), .S0(n65872), 
        .S1(n65766), .Q(n30875) );
  IMUX40 U70221 ( .A(n65628), .B(n65629), .C(n65630), .D(n65631), .S0(n65890), 
        .S1(n65747), .Q(n63505) );
  IMUX40 U70217 ( .A(n65612), .B(n65613), .C(n65614), .D(n65615), .S0(n65854), 
        .S1(n65753), .Q(n63500) );
  IMUX40 U71565 ( .A(n65628), .B(n65629), .C(n65630), .D(n65631), .S0(n65890), 
        .S1(n65766), .Q(n64785) );
  IMUX40 U71561 ( .A(n65612), .B(n65613), .C(n65614), .D(n65615), .S0(n65876), 
        .S1(n65765), .Q(n64780) );
  IMUX40 U68205 ( .A(n65628), .B(n65629), .C(n65630), .D(n65631), .S0(n65902), 
        .S1(n65766), .Q(n61585) );
  IMUX40 U68201 ( .A(n65612), .B(n65613), .C(n65614), .D(n65615), .S0(n65877), 
        .S1(n65770), .Q(n61580) );
  IMUX40 U68213 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65848), 
        .S1(n65762), .Q(n61595) );
  IMUX40 U70893 ( .A(n65628), .B(n65629), .C(n65630), .D(n65631), .S0(n65795), 
        .S1(N1256), .Q(n64145) );
  IMUX40 U70889 ( .A(n65612), .B(n65613), .C(n65614), .D(n65615), .S0(n65810), 
        .S1(N1256), .Q(n64140) );
  IMUX40 U70901 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65801), 
        .S1(N1256), .Q(n64155) );
  IMUX40 U37293 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(n65783), 
        .S1(N956), .Q(n32145) );
  IMUX40 U37289 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65803), 
        .S1(N956), .Q(n32140) );
  IMUX40 U37297 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65797), 
        .S1(N956), .Q(n32150) );
  IMUX40 U69549 ( .A(n65628), .B(n65629), .C(n65630), .D(n65631), .S0(n65825), 
        .S1(N1244), .Q(n62865) );
  IMUX40 U69553 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65813), 
        .S1(N1244), .Q(n62870) );
  IMUX40 U38637 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(n65782), 
        .S1(N968), .Q(n33425) );
  IMUX40 U38633 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65816), 
        .S1(N968), .Q(n33420) );
  IMUX40 U38645 ( .A(n65724), .B(n65725), .C(n65726), .D(n65727), .S0(n65822), 
        .S1(N968), .Q(n33435) );
  IMUX40 U69545 ( .A(n65612), .B(n65613), .C(n65614), .D(n65615), .S0(n65805), 
        .S1(N1244), .Q(n62860) );
  IMUX40 U37964 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65877), 
        .S1(n65745), .Q(n32787) );
  IMUX40 U37960 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65878), 
        .S1(n65756), .Q(n32782) );
  IMUX40 U37972 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65904), 
        .S1(n65753), .Q(n32797) );
  IMUX40 U37968 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65905), 
        .S1(n65744), .Q(n32792) );
  IMUX40 U39308 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65904), 
        .S1(n65768), .Q(n34067) );
  IMUX40 U39304 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65885), 
        .S1(n65767), .Q(n34062) );
  IMUX40 U39316 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65874), 
        .S1(n65769), .Q(n34077) );
  IMUX40 U39312 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65845), 
        .S1(n65769), .Q(n34072) );
  IMUX40 U36620 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65888), 
        .S1(n65755), .Q(n31507) );
  IMUX40 U36616 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65845), 
        .S1(n65755), .Q(n31502) );
  IMUX40 U36628 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65869), 
        .S1(n65756), .Q(n31517) );
  IMUX40 U36624 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65884), 
        .S1(n65756), .Q(n31512) );
  IMUX40 U35948 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65873), 
        .S1(n65768), .Q(n30867) );
  IMUX40 U35944 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65874), 
        .S1(n65760), .Q(n30862) );
  IMUX40 U35956 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65872), 
        .S1(n65772), .Q(n30877) );
  IMUX40 U35952 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65858), 
        .S1(n65761), .Q(n30872) );
  IMUX40 U70220 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65895), 
        .S1(n65753), .Q(n63507) );
  IMUX40 U70216 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65879), 
        .S1(n65753), .Q(n63502) );
  IMUX40 U70228 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65850), 
        .S1(n65748), .Q(n63517) );
  IMUX40 U70224 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65851), 
        .S1(n65757), .Q(n63512) );
  IMUX40 U71564 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65854), 
        .S1(n65765), .Q(n64787) );
  IMUX40 U71560 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65866), 
        .S1(n65765), .Q(n64782) );
  IMUX40 U71572 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65895), 
        .S1(n65767), .Q(n64797) );
  IMUX40 U71568 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65906), 
        .S1(n65766), .Q(n64792) );
  IMUX40 U68876 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65894), 
        .S1(n65757), .Q(n62227) );
  IMUX40 U68872 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65900), 
        .S1(n65756), .Q(n62222) );
  IMUX40 U68884 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65879), 
        .S1(n65757), .Q(n62237) );
  IMUX40 U68880 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65889), 
        .S1(n65757), .Q(n62232) );
  IMUX40 U68204 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65866), 
        .S1(n65761), .Q(n61587) );
  IMUX40 U68200 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65851), 
        .S1(n65762), .Q(n61582) );
  IMUX40 U68212 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65832), 
        .S1(n65769), .Q(n61597) );
  IMUX40 U68208 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65848), 
        .S1(n65775), .Q(n61592) );
  IMUX40 U49389 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65835), .S1(n65745), .Q(n43665) );
  IMUX40 U49385 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65891), .S1(n65755), .Q(n43660) );
  IMUX40 U49397 ( .A(\OFill[0][0] ), .B(n65661), .C(n65662), .D(n65663), .S0(
        n65895), .S1(n65754), .Q(n43675) );
  IMUX40 U50061 ( .A(n65628), .B(n65629), .C(n65630), .D(n65631), .S0(n65841), 
        .S1(n65756), .Q(n44305) );
  IMUX40 U50057 ( .A(\OFill[48][0] ), .B(n65613), .C(n65614), .D(n65615), .S0(
        n65840), .S1(n65754), .Q(n44300) );
  IMUX40 U50069 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65844), .S1(n65753), .Q(n44315) );
  IMUX40 U51405 ( .A(n65628), .B(\OFill[33][0] ), .C(\OFill[34][0] ), .D(
        \OFill[35][0] ), .S0(n65813), .S1(n65922), .Q(n45585) );
  IMUX40 U51401 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65818), .S1(n65538), .Q(n45580) );
  IMUX40 U51413 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65795), 
        .S1(n65922), .Q(n45595) );
  IMUX40 U62829 ( .A(n65628), .B(n65629), .C(\OFill[34][0] ), .D(n65631), .S0(
        n65786), .S1(N1184), .Q(n56465) );
  IMUX40 U62825 ( .A(n65612), .B(n65613), .C(\OFill[50][0] ), .D(n65615), .S0(
        n65788), .S1(n65913), .Q(n56460) );
  IMUX40 U62837 ( .A(n65660), .B(\OFill[1][0] ), .C(n65662), .D(n65663), .S0(
        n65805), .S1(N968), .Q(n56475) );
  IMUX40 U62157 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65867), .S1(N1208), .Q(n55825) );
  IMUX40 U62153 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65876), .S1(n65746), .Q(n55820) );
  IMUX40 U62165 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65896), .S1(n65745), .Q(n55835) );
  IMUX40 U63501 ( .A(n65628), .B(n65629), .C(\OFill[34][0] ), .D(n65631), .S0(
        n65841), .S1(n65764), .Q(n57105) );
  IMUX40 U63497 ( .A(n65612), .B(n65613), .C(\OFill[50][0] ), .D(n65615), .S0(
        n65898), .S1(n65772), .Q(n57100) );
  IMUX40 U63509 ( .A(n65660), .B(\OFill[1][0] ), .C(n65662), .D(n65663), .S0(
        n65856), .S1(n65761), .Q(n57115) );
  IMUX40 U64173 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65851), .S1(n65764), .Q(n57745) );
  IMUX40 U64169 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65845), .S1(n65768), .Q(n57740) );
  IMUX40 U64181 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65894), .S1(n65776), .Q(n57755) );
  IMUX40 U65517 ( .A(n65628), .B(n65629), .C(\OFill[34][0] ), .D(
        \OFill[35][0] ), .S0(n65856), .S1(n65750), .Q(n59025) );
  IMUX40 U65513 ( .A(n65612), .B(n65613), .C(\OFill[50][0] ), .D(
        \OFill[51][0] ), .S0(n65894), .S1(n65753), .Q(n59020) );
  IMUX40 U65525 ( .A(n65660), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65879), .S1(n65749), .Q(n59035) );
  IMUX40 U17133 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65857), .S1(n65756), .Q(n12945) );
  IMUX40 U17129 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65878), .S1(n65744), .Q(n12940) );
  IMUX40 U17141 ( .A(\GFill[0][0] ), .B(n65725), .C(n65726), .D(n65727), .S0(
        n65902), .S1(n65757), .Q(n12955) );
  IMUX40 U16461 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(n65786), 
        .S1(n65911), .Q(n12305) );
  IMUX40 U16457 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65788), 
        .S1(n65912), .Q(n12300) );
  IMUX40 U16469 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65814), .S1(n65912), .Q(n12315) );
  IMUX40 U18477 ( .A(n65692), .B(\GFill[33][0] ), .C(\GFill[34][0] ), .D(
        \GFill[35][0] ), .S0(N1207), .S1(n65768), .Q(n14225) );
  IMUX40 U18473 ( .A(n65676), .B(\GFill[49][0] ), .C(\GFill[50][0] ), .D(
        \GFill[51][0] ), .S0(n65891), .S1(n65770), .Q(n14220) );
  IMUX40 U18485 ( .A(n65724), .B(n65725), .C(n65726), .D(n65727), .S0(n65889), 
        .S1(n65771), .Q(n14235) );
  IMUX40 U17805 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(n65695), .S0(n65836), .S1(n65753), .Q(n13585) );
  IMUX40 U17801 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(n65679), .S0(n65837), .S1(n65752), .Q(n13580) );
  IMUX40 U17813 ( .A(n65724), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65833), .S1(n65746), .Q(n13595) );
  IMUX40 U19149 ( .A(n65692), .B(n65693), .C(n65694), .D(\GFill[35][0] ), .S0(
        n65793), .S1(N1082), .Q(n14865) );
  IMUX40 U19145 ( .A(n65676), .B(n65677), .C(n65678), .D(\GFill[51][0] ), .S0(
        n65797), .S1(n65743), .Q(n14860) );
  IMUX40 U19157 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        n65727), .S0(n65804), .S1(n65912), .Q(n14875) );
  IMUX40 U30573 ( .A(n65692), .B(\GFill[33][0] ), .C(n65694), .D(
        \GFill[35][0] ), .S0(n65817), .S1(n65921), .Q(n25745) );
  IMUX40 U30569 ( .A(n65676), .B(\GFill[49][0] ), .C(n65678), .D(
        \GFill[51][0] ), .S0(n65826), .S1(n65913), .Q(n25740) );
  IMUX40 U30581 ( .A(n65724), .B(n65725), .C(\GFill[2][0] ), .D(n65727), .S0(
        n65787), .S1(N1112), .Q(n25755) );
  IMUX40 U29901 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65838), .S1(n65752), .Q(n25105) );
  IMUX40 U29897 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65846), .S1(n65752), .Q(n25100) );
  IMUX40 U29909 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65888), .S1(n65756), .Q(n25115) );
  IMUX40 U31245 ( .A(n65692), .B(\GFill[33][0] ), .C(n65694), .D(
        \GFill[35][0] ), .S0(n65876), .S1(n65762), .Q(n26385) );
  IMUX40 U31241 ( .A(n65676), .B(\GFill[49][0] ), .C(n65678), .D(
        \GFill[51][0] ), .S0(n65858), .S1(n65768), .Q(n26380) );
  IMUX40 U31253 ( .A(n65724), .B(n65725), .C(\GFill[2][0] ), .D(n65727), .S0(
        n65893), .S1(n65777), .Q(n26395) );
  IMUX40 U32589 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65814), .S1(n65534), .Q(n27665) );
  IMUX40 U32585 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65788), .S1(n65538), .Q(n27660) );
  IMUX40 U32597 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65806), .S1(N1148), .Q(n27675) );
  IMUX40 U31917 ( .A(n65692), .B(\GFill[33][0] ), .C(n65694), .D(
        \GFill[35][0] ), .S0(n65860), .S1(n65778), .Q(n27025) );
  IMUX40 U31913 ( .A(n65676), .B(\GFill[49][0] ), .C(n65678), .D(
        \GFill[51][0] ), .S0(n65909), .S1(n65772), .Q(n27020) );
  IMUX40 U31925 ( .A(n65724), .B(n65725), .C(\GFill[2][0] ), .D(\GFill[3][0] ), 
        .S0(n65908), .S1(n65771), .Q(n27035) );
  IMUX40 U33261 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65890), .S1(n65752), .Q(n28305) );
  IMUX40 U33257 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65886), .S1(n65747), .Q(n28300) );
  IMUX40 U33269 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        n65727), .S0(n65855), .S1(n65744), .Q(n28315) );
  IMUX40 U23181 ( .A(\GFill[32][0] ), .B(n65693), .C(n65694), .D(
        \GFill[35][0] ), .S0(n65909), .S1(n65751), .Q(n18705) );
  IMUX40 U23177 ( .A(\GFill[48][0] ), .B(n65677), .C(n65678), .D(
        \GFill[51][0] ), .S0(n65862), .S1(n65750), .Q(n18700) );
  IMUX40 U23189 ( .A(n65724), .B(n65725), .C(n65726), .D(\GFill[3][0] ), .S0(
        n65896), .S1(n65756), .Q(n18715) );
  IMUX40 U22509 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65792), .S1(n65913), .Q(n18065) );
  IMUX40 U22505 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65803), .S1(N1184), .Q(n18060) );
  IMUX40 U22517 ( .A(\GFill[0][0] ), .B(n65725), .C(n65726), .D(\GFill[3][0] ), 
        .S0(n65816), .S1(N1184), .Q(n18075) );
  IMUX40 U35277 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(n65835), 
        .S1(n65754), .Q(n30225) );
  IMUX40 U35273 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65880), 
        .S1(n65754), .Q(n30220) );
  IMUX40 U54093 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(n65631), .S0(n65852), .S1(n65772), .Q(n48145) );
  IMUX40 U54089 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(n65615), .S0(n65851), .S1(n65769), .Q(n48140) );
  IMUX40 U54101 ( .A(n65660), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65854), .S1(n65773), .Q(n48155) );
  IMUX40 U55437 ( .A(n65628), .B(n65629), .C(n65630), .D(\OFill[35][0] ), .S0(
        n65885), .S1(n65754), .Q(n49425) );
  IMUX40 U55433 ( .A(\OFill[48][0] ), .B(n65613), .C(n65614), .D(
        \OFill[51][0] ), .S0(n65839), .S1(n65756), .Q(n49420) );
  IMUX40 U55445 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(n65662), .D(n65663), 
        .S0(n65851), .S1(n65749), .Q(n49435) );
  IMUX40 U67533 ( .A(\OFill[32][0] ), .B(n65629), .C(n65630), .D(n65631), .S0(
        n65899), .S1(n65747), .Q(n60945) );
  IMUX40 U67529 ( .A(\OFill[48][0] ), .B(n65613), .C(n65614), .D(n65615), .S0(
        n65871), .S1(n65747), .Q(n60940) );
  IMUX40 U9069 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65811), .S1(N704), .Q(n5265) );
  IMUX40 U9065 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65808), .S1(N704), .Q(n5260) );
  IMUX40 U8397 ( .A(\GFill[32][0] ), .B(n65693), .C(\GFill[34][0] ), .D(n65695), .S0(n65809), .S1(n65536), .Q(n4625) );
  IMUX40 U8393 ( .A(\GFill[48][0] ), .B(n65677), .C(\GFill[50][0] ), .D(n65679), .S0(n65810), .S1(n65536), .Q(n4620) );
  IMUX40 U8405 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(n65726), .D(
        \GFill[3][0] ), .S0(n65789), .S1(n65536), .Q(n4635) );
  IMUX40 U10413 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65818), .S1(N716), .Q(n6545) );
  IMUX40 U10409 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65819), .S1(N716), .Q(n6540) );
  IMUX40 U9741 ( .A(\GFill[32][0] ), .B(n65693), .C(\GFill[34][0] ), .D(
        \GFill[35][0] ), .S0(n65800), .S1(n65935), .Q(n5905) );
  IMUX40 U9737 ( .A(\GFill[48][0] ), .B(n65677), .C(\GFill[50][0] ), .D(
        \GFill[51][0] ), .S0(n65799), .S1(n65934), .Q(n5900) );
  IMUX40 U9749 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65798), .S1(n65935), .Q(n5915) );
  IMUX40 U11085 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(n65695), .S0(n65831), .S1(N722), .Q(n7185) );
  IMUX40 U11081 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(n65679), .S0(n65829), .S1(N722), .Q(n7180) );
  IMUX40 U12429 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(n65695), .S0(n65805), .S1(N1016), .Q(n8465) );
  IMUX40 U12425 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(n65679), .S0(n65804), .S1(n65930), .Q(n8460) );
  IMUX40 U12437 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(n65726), .D(
        \GFill[3][0] ), .S0(n65803), .S1(n65933), .Q(n8475) );
  IMUX40 U11757 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65822), .S1(n65932), .Q(n7825) );
  IMUX40 U11753 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65829), .S1(n65931), .Q(n7820) );
  IMUX40 U11765 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65795), .S1(n65931), .Q(n7835) );
  IMUX40 U13773 ( .A(n65692), .B(\GFill[33][0] ), .C(\GFill[34][0] ), .D(
        n65695), .S0(n65792), .S1(n65929), .Q(n9745) );
  IMUX40 U13769 ( .A(n65676), .B(\GFill[49][0] ), .C(\GFill[50][0] ), .D(
        n65679), .S0(n65791), .S1(n65928), .Q(n9740) );
  IMUX40 U13781 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(n65726), .D(
        \GFill[3][0] ), .S0(n65790), .S1(n65929), .Q(n9755) );
  IMUX40 U15117 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65796), .S1(N1010), .Q(n11025) );
  IMUX40 U15113 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65796), .S1(n65925), .Q(n11020) );
  IMUX40 U15125 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65795), .S1(N1046), .Q(n11035) );
  IMUX40 U14445 ( .A(n65692), .B(\GFill[33][0] ), .C(n65694), .D(
        \GFill[35][0] ), .S0(n65807), .S1(n65927), .Q(n10385) );
  IMUX40 U14441 ( .A(n65676), .B(\GFill[49][0] ), .C(n65678), .D(
        \GFill[51][0] ), .S0(n65807), .S1(n65926), .Q(n10380) );
  IMUX40 U14453 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65813), .S1(n65927), .Q(n10395) );
  IMUX40 U27885 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65891), .S1(n65772), .Q(n23185) );
  IMUX40 U27881 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65897), .S1(n65772), .Q(n23180) );
  IMUX40 U29229 ( .A(n65692), .B(\GFill[33][0] ), .C(\GFill[34][0] ), .D(
        \GFill[35][0] ), .S0(n65796), .S1(N1112), .Q(n24465) );
  IMUX40 U29225 ( .A(n65676), .B(\GFill[49][0] ), .C(\GFill[50][0] ), .D(
        \GFill[51][0] ), .S0(n65782), .S1(N1244), .Q(n24460) );
  IMUX40 U29237 ( .A(n65724), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(n65727), 
        .S0(n65802), .S1(N1112), .Q(n24475) );
  IMUX40 U25869 ( .A(n65692), .B(\GFill[33][0] ), .C(\GFill[34][0] ), .D(
        n65695), .S0(n65910), .S1(n65779), .Q(n21265) );
  IMUX40 U25865 ( .A(n65676), .B(\GFill[49][0] ), .C(\GFill[50][0] ), .D(
        n65679), .S0(n65833), .S1(n65765), .Q(n21260) );
  IMUX40 U27213 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65835), .S1(n65746), .Q(n22545) );
  IMUX40 U27209 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65863), .S1(n65745), .Q(n22540) );
  IMUX40 U27221 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65910), .S1(n65746), .Q(n22555) );
  IMUX40 U24525 ( .A(\GFill[32][0] ), .B(n65693), .C(n65694), .D(
        \GFill[35][0] ), .S0(n65804), .S1(N842), .Q(n19985) );
  IMUX40 U24521 ( .A(\GFill[48][0] ), .B(n65677), .C(n65678), .D(
        \GFill[51][0] ), .S0(n65814), .S1(N842), .Q(n19980) );
  IMUX40 U24533 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65785), .S1(N842), .Q(n19995) );
  IMUX40 U23853 ( .A(n65692), .B(\GFill[33][0] ), .C(\GFill[34][0] ), .D(
        \GFill[35][0] ), .S0(n65861), .S1(n65763), .Q(n19345) );
  IMUX40 U23849 ( .A(n65676), .B(\GFill[49][0] ), .C(\GFill[50][0] ), .D(
        \GFill[51][0] ), .S0(n65847), .S1(n65778), .Q(n19340) );
  IMUX40 U23861 ( .A(n65724), .B(n65725), .C(n65726), .D(\GFill[3][0] ), .S0(
        n65889), .S1(n65766), .Q(n19355) );
  IMUX40 U41325 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(n65630), .D(
        \OFill[35][0] ), .S0(n65816), .S1(N1004), .Q(n35985) );
  IMUX40 U41321 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(n65614), .D(
        \OFill[51][0] ), .S0(n65817), .S1(N1004), .Q(n35980) );
  IMUX40 U42669 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65828), .S1(N1034), .Q(n37265) );
  IMUX40 U42665 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65828), .S1(N1034), .Q(n37260) );
  IMUX40 U41997 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(n65630), .D(
        \OFill[35][0] ), .S0(n65801), .S1(n65935), .Q(n36625) );
  IMUX40 U41993 ( .A(n65612), .B(\OFill[49][0] ), .C(n65614), .D(
        \OFill[51][0] ), .S0(n65798), .S1(n65934), .Q(n36620) );
  IMUX40 U42005 ( .A(\OFill[0][0] ), .B(n65661), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65800), .S1(n65934), .Q(n36635) );
  IMUX40 U43341 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65826), .S1(N1010), .Q(n37905) );
  IMUX40 U43337 ( .A(n65612), .B(\OFill[49][0] ), .C(\OFill[50][0] ), .D(
        \OFill[51][0] ), .S0(n65825), .S1(N980), .Q(n37900) );
  IMUX40 U44685 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(n65630), .D(
        \OFill[35][0] ), .S0(n65806), .S1(n65932), .Q(n39185) );
  IMUX40 U44681 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(n65614), .D(
        \OFill[51][0] ), .S0(n65803), .S1(n65933), .Q(n39180) );
  IMUX40 U44693 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65805), .S1(n65930), .Q(n39195) );
  IMUX40 U44013 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65816), .S1(n65933), .Q(n38545) );
  IMUX40 U44009 ( .A(n65612), .B(\OFill[49][0] ), .C(\OFill[50][0] ), .D(
        \OFill[51][0] ), .S0(n65797), .S1(n65930), .Q(n38540) );
  IMUX40 U44021 ( .A(\OFill[0][0] ), .B(n65661), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65806), .S1(n65931), .Q(n38555) );
  IMUX40 U45357 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65821), .S1(N1040), .Q(n39825) );
  IMUX40 U45353 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65821), .S1(N1040), .Q(n39820) );
  IMUX40 U46701 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65782), .S1(n65927), .Q(n41105) );
  IMUX40 U46697 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65812), .S1(n65926), .Q(n41100) );
  IMUX40 U46709 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65829), .S1(n65926), .Q(n41115) );
  IMUX40 U46029 ( .A(n65628), .B(\OFill[33][0] ), .C(\OFill[34][0] ), .D(
        n65631), .S0(n65793), .S1(n65929), .Q(n40465) );
  IMUX40 U46025 ( .A(n65612), .B(\OFill[49][0] ), .C(\OFill[50][0] ), .D(
        n65615), .S0(n65790), .S1(n65928), .Q(n40460) );
  IMUX40 U46037 ( .A(\OFill[0][0] ), .B(n65661), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65792), .S1(n65928), .Q(n40475) );
  IMUX40 U47373 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65813), .S1(N1010), .Q(n41745) );
  IMUX40 U47369 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65795), .S1(n65925), .Q(n41740) );
  IMUX40 U47381 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65796), .S1(n65924), .Q(n41755) );
  IMUX40 U60141 ( .A(n65628), .B(\OFill[33][0] ), .C(\OFill[34][0] ), .D(
        n65631), .S0(N1207), .S1(n65771), .Q(n53905) );
  IMUX40 U60137 ( .A(n65612), .B(\OFill[49][0] ), .C(\OFill[50][0] ), .D(
        n65615), .S0(n65906), .S1(n65770), .Q(n53900) );
  IMUX40 U61485 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(n65631), .S0(n65826), .S1(N1112), .Q(n55185) );
  IMUX40 U61481 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(n65615), .S0(n65825), .S1(n65913), .Q(n55180) );
  IMUX40 U61493 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(n65662), .D(n65663), 
        .S0(n65817), .S1(N956), .Q(n55195) );
  IMUX40 U58125 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65892), .S1(n65773), .Q(n51985) );
  IMUX40 U58121 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65877), .S1(n65773), .Q(n51980) );
  IMUX40 U59469 ( .A(n65628), .B(\OFill[33][0] ), .C(\OFill[34][0] ), .D(
        n65631), .S0(n65844), .S1(n65745), .Q(n53265) );
  IMUX40 U59465 ( .A(n65612), .B(\OFill[49][0] ), .C(\OFill[50][0] ), .D(
        n65615), .S0(n65895), .S1(n65745), .Q(n53260) );
  IMUX40 U59477 ( .A(n65660), .B(\OFill[1][0] ), .C(n65662), .D(n65663), .S0(
        n65900), .S1(n65744), .Q(n53275) );
  IMUX40 U56109 ( .A(\OFill[32][0] ), .B(n65629), .C(n65630), .D(
        \OFill[35][0] ), .S0(n65876), .S1(n65763), .Q(n50065) );
  IMUX40 U56105 ( .A(\OFill[48][0] ), .B(n65613), .C(n65614), .D(
        \OFill[51][0] ), .S0(n65859), .S1(n65772), .Q(n50060) );
  IMUX40 U57453 ( .A(n65628), .B(\OFill[33][0] ), .C(\OFill[34][0] ), .D(
        \OFill[35][0] ), .S0(n65891), .S1(n65748), .Q(n51345) );
  IMUX40 U57449 ( .A(n65612), .B(\OFill[49][0] ), .C(\OFill[50][0] ), .D(
        \OFill[51][0] ), .S0(n65882), .S1(n65748), .Q(n51340) );
  IMUX40 U23185 ( .A(\GFill[16][0] ), .B(n65709), .C(n65710), .D(n65711), .S0(
        n65852), .S1(n65747), .Q(n18710) );
  IMUX40 U23182 ( .A(\GFill[28][0] ), .B(n65721), .C(n65722), .D(n65723), .S0(
        n65883), .S1(n65751), .Q(n18713) );
  IMUX40 U23183 ( .A(\GFill[24][0] ), .B(n65717), .C(n65718), .D(n65719), .S0(
        n65842), .S1(N1208), .Q(n18711) );
  IMUX40 U23016 ( .A(n18710), .B(n18711), .C(n18712), .D(n18713), .S0(N1120), 
        .S1(n65917), .Q(n18709) );
  IMUX40 U55441 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65864), 
        .S1(n65749), .Q(n49430) );
  IMUX40 U55438 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65885), 
        .S1(n65749), .Q(n49433) );
  IMUX40 U55439 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65896), 
        .S1(n65749), .Q(n49431) );
  IMUX40 U55272 ( .A(n49430), .B(n49431), .C(n49432), .D(n49433), .S0(N11412), 
        .S1(n65917), .Q(n49429) );
  IMUX40 U23857 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65903), .S1(n65761), .Q(n19350) );
  IMUX40 U23854 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65908), .S1(n65778), .Q(n19353) );
  IMUX40 U23855 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65887), .S1(n65781), .Q(n19351) );
  IMUX40 U23688 ( .A(n19350), .B(n19351), .C(n19352), .D(n19353), .S0(N838), 
        .S1(N837), .Q(n19349) );
  IMUX40 U25205 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65878), .S1(n65754), .Q(n20635) );
  IMUX40 U25202 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65857), .S1(n65753), .Q(n20638) );
  IMUX40 U25203 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65861), .S1(n65754), .Q(n20636) );
  IMUX40 U25033 ( .A(n20635), .B(n20636), .C(n20637), .D(n20638), .S0(N850), 
        .S1(n65919), .Q(n20634) );
  IMUX40 U25201 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65898), 
        .S1(n65753), .Q(n20630) );
  IMUX40 U25198 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65856), 
        .S1(n65753), .Q(n20633) );
  IMUX40 U25199 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65856), 
        .S1(n65753), .Q(n20631) );
  IMUX40 U25032 ( .A(n20630), .B(n20631), .C(n20632), .D(n20633), .S0(N850), 
        .S1(n65919), .Q(n20629) );
  IMUX40 U70892 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65788), 
        .S1(N1256), .Q(n64147) );
  IMUX40 U70888 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65800), 
        .S1(N1256), .Q(n64142) );
  IMUX40 U70900 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65808), 
        .S1(N1256), .Q(n64157) );
  IMUX40 U70896 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65809), 
        .S1(N1256), .Q(n64152) );
  IMUX40 U37292 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65816), 
        .S1(N956), .Q(n32147) );
  IMUX40 U37288 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65827), 
        .S1(N956), .Q(n32142) );
  IMUX40 U37296 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65796), 
        .S1(N956), .Q(n32152) );
  IMUX40 U37300 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65794), 
        .S1(N956), .Q(n32157) );
  IMUX40 U69548 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65804), 
        .S1(N1244), .Q(n62867) );
  IMUX40 U69552 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65828), 
        .S1(N1244), .Q(n62872) );
  IMUX40 U38636 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65787), 
        .S1(N968), .Q(n33427) );
  IMUX40 U38632 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65798), 
        .S1(N968), .Q(n33422) );
  IMUX40 U38644 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65786), 
        .S1(N968), .Q(n33437) );
  IMUX40 U38640 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65830), 
        .S1(N968), .Q(n33432) );
  IMUX40 U69544 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65783), 
        .S1(N1244), .Q(n62862) );
  IMUX40 U69556 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65818), 
        .S1(N1244), .Q(n62877) );
  IMUX40 U48716 ( .A(\OFill[36][0] ), .B(n65633), .C(n65634), .D(n65635), .S0(
        n65819), .S1(n65743), .Q(n43027) );
  IMUX40 U48712 ( .A(\OFill[52][0] ), .B(n65617), .C(n65618), .D(n65619), .S0(
        n65804), .S1(N1220), .Q(n43022) );
  IMUX40 U48724 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65783), 
        .S1(n65911), .Q(n43037) );
  IMUX40 U48720 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65826), 
        .S1(n65912), .Q(n43032) );
  IMUX40 U48044 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65866), .S1(n65778), .Q(n42387) );
  IMUX40 U48040 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65865), .S1(n65777), .Q(n42382) );
  IMUX40 U48052 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65833), .S1(n65761), .Q(n42397) );
  IMUX40 U48048 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65852), .S1(n65776), .Q(n42392) );
  IMUX40 U49388 ( .A(\OFill[36][0] ), .B(n65633), .C(n65634), .D(n65635), .S0(
        n65901), .S1(N1208), .Q(n43667) );
  IMUX40 U49384 ( .A(\OFill[52][0] ), .B(n65617), .C(n65618), .D(n65619), .S0(
        n65882), .S1(n65753), .Q(n43662) );
  IMUX40 U49396 ( .A(\OFill[4][0] ), .B(n65665), .C(n65666), .D(n65667), .S0(
        n65876), .S1(N1208), .Q(n43677) );
  IMUX40 U49392 ( .A(\OFill[20][0] ), .B(n65649), .C(n65650), .D(n65651), .S0(
        n65910), .S1(N1208), .Q(n43672) );
  IMUX40 U50732 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65885), .S1(n65762), .Q(n44947) );
  IMUX40 U50728 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65872), .S1(n65770), .Q(n44942) );
  IMUX40 U50740 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65879), .S1(n65772), .Q(n44957) );
  IMUX40 U50736 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65891), .S1(n65779), .Q(n44952) );
  IMUX40 U50060 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(n65635), .S0(n65841), .S1(n65747), .Q(n44307) );
  IMUX40 U50056 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(n65619), .S0(n65839), .S1(n65752), .Q(n44302) );
  IMUX40 U50068 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(n65666), .D(n65667), 
        .S0(n65843), .S1(n65748), .Q(n44317) );
  IMUX40 U50064 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65842), .S1(n65744), .Q(n44312) );
  IMUX40 U51404 ( .A(\OFill[36][0] ), .B(n65633), .C(n65634), .D(
        \OFill[39][0] ), .S0(n65812), .S1(n65922), .Q(n45587) );
  IMUX40 U51400 ( .A(\OFill[52][0] ), .B(n65617), .C(n65618), .D(
        \OFill[55][0] ), .S0(n65817), .S1(n65912), .Q(n45582) );
  IMUX40 U51412 ( .A(n65664), .B(n65665), .C(\OFill[6][0] ), .D(\OFill[7][0] ), 
        .S0(n65796), .S1(n65922), .Q(n45597) );
  IMUX40 U51408 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(n65820), 
        .S1(n65922), .Q(n45592) );
  IMUX40 U62828 ( .A(n65632), .B(n65633), .C(\OFill[38][0] ), .D(n65635), .S0(
        n65789), .S1(n65921), .Q(n56467) );
  IMUX40 U62824 ( .A(n65616), .B(n65617), .C(\OFill[54][0] ), .D(n65619), .S0(
        n65825), .S1(n65921), .Q(n56462) );
  IMUX40 U62836 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(n65666), .D(n65667), 
        .S0(n65800), .S1(N1112), .Q(n56477) );
  IMUX40 U62832 ( .A(\OFill[20][0] ), .B(n65649), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65803), .S1(N1172), .Q(n56472) );
  IMUX40 U62156 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65873), .S1(n65744), .Q(n55827) );
  IMUX40 U62152 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65903), .S1(n65752), .Q(n55822) );
  IMUX40 U62164 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65869), .S1(n65749), .Q(n55837) );
  IMUX40 U62160 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65868), .S1(n65751), .Q(n55832) );
  IMUX40 U63500 ( .A(n65632), .B(n65633), .C(\OFill[38][0] ), .D(n65635), .S0(
        n65837), .S1(n65769), .Q(n57107) );
  IMUX40 U63496 ( .A(n65616), .B(n65617), .C(\OFill[54][0] ), .D(n65619), .S0(
        n65848), .S1(n65759), .Q(n57102) );
  IMUX40 U63508 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(n65666), .D(n65667), 
        .S0(n65895), .S1(n65767), .Q(n57117) );
  IMUX40 U63504 ( .A(n65648), .B(n65649), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65860), .S1(n65770), .Q(n57112) );
  IMUX40 U64844 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65804), .S1(N1082), .Q(n58387) );
  IMUX40 U64840 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65828), .S1(n65743), .Q(n58382) );
  IMUX40 U64852 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65790), .S1(n65911), .Q(n58397) );
  IMUX40 U64848 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65804), .S1(n65911), .Q(n58392) );
  IMUX40 U64172 ( .A(n65632), .B(n65633), .C(\OFill[38][0] ), .D(
        \OFill[39][0] ), .S0(n65898), .S1(n65767), .Q(n57747) );
  IMUX40 U64168 ( .A(n65616), .B(n65617), .C(\OFill[54][0] ), .D(
        \OFill[55][0] ), .S0(n65908), .S1(n65766), .Q(n57742) );
  IMUX40 U64180 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65901), .S1(n65772), .Q(n57757) );
  IMUX40 U64176 ( .A(\OFill[20][0] ), .B(n65649), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65859), .S1(n65777), .Q(n57752) );
  IMUX40 U65516 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(n65635), .S0(n65863), .S1(N1208), .Q(n59027) );
  IMUX40 U65512 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(n65619), .S0(n65856), .S1(n65748), .Q(n59022) );
  IMUX40 U65524 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(n65666), .D(n65667), 
        .S0(N1207), .S1(N1208), .Q(n59037) );
  IMUX40 U65520 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65905), .S1(n65757), .Q(n59032) );
  IMUX40 U15788 ( .A(\GFill[36][0] ), .B(n65697), .C(n65698), .D(n65699), .S0(
        n65862), .S1(n65767), .Q(n11667) );
  IMUX40 U15784 ( .A(\GFill[52][0] ), .B(n65681), .C(n65682), .D(n65683), .S0(
        n65863), .S1(n65768), .Q(n11662) );
  IMUX40 U15796 ( .A(\GFill[4][0] ), .B(n65729), .C(\GFill[6][0] ), .D(n65731), 
        .S0(n65859), .S1(n65774), .Q(n11677) );
  IMUX40 U15792 ( .A(\GFill[20][0] ), .B(n65713), .C(n65714), .D(n65715), .S0(
        n65860), .S1(n65762), .Q(n11672) );
  IMUX40 U17132 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65901), .S1(n65753), .Q(n12947) );
  IMUX40 U17128 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65908), .S1(n65756), .Q(n12942) );
  IMUX40 U17140 ( .A(n65728), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65892), .S1(n65747), .Q(n12957) );
  IMUX40 U17136 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65858), .S1(n65748), .Q(n12952) );
  IMUX40 U16460 ( .A(\GFill[36][0] ), .B(n65697), .C(n65698), .D(n65699), .S0(
        n65786), .S1(n65743), .Q(n12307) );
  IMUX40 U16456 ( .A(\GFill[52][0] ), .B(n65681), .C(n65682), .D(n65683), .S0(
        n65785), .S1(N1082), .Q(n12302) );
  IMUX40 U16468 ( .A(\GFill[4][0] ), .B(n65729), .C(\GFill[6][0] ), .D(n65731), 
        .S0(n65815), .S1(n65912), .Q(n12317) );
  IMUX40 U16464 ( .A(\GFill[20][0] ), .B(n65713), .C(n65714), .D(n65715), .S0(
        n65813), .S1(N1082), .Q(n12312) );
  IMUX40 U18476 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65900), .S1(n65774), .Q(n14227) );
  IMUX40 U18472 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65848), .S1(n65773), .Q(n14222) );
  IMUX40 U18484 ( .A(n65728), .B(n65729), .C(\GFill[6][0] ), .D(\GFill[7][0] ), 
        .S0(N1207), .S1(n65781), .Q(n14237) );
  IMUX40 U18480 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65910), .S1(n65778), .Q(n14232) );
  IMUX40 U17804 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(n65699), .S0(n65836), .S1(n65749), .Q(n13587) );
  IMUX40 U17800 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(n65683), .S0(n65838), .S1(n65751), .Q(n13582) );
  IMUX40 U17812 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        n65731), .S0(n65834), .S1(n65744), .Q(n13597) );
  IMUX40 U17808 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(n65715), .S0(n65835), .S1(n65746), .Q(n13592) );
  IMUX40 U19148 ( .A(\GFill[36][0] ), .B(n65697), .C(n65698), .D(
        \GFill[39][0] ), .S0(n65826), .S1(n65538), .Q(n14867) );
  IMUX40 U19144 ( .A(\GFill[52][0] ), .B(n65681), .C(n65682), .D(
        \GFill[55][0] ), .S0(n65819), .S1(n65923), .Q(n14862) );
  IMUX40 U19156 ( .A(n65728), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65810), .S1(n65743), .Q(n14877) );
  IMUX40 U19152 ( .A(\GFill[20][0] ), .B(n65713), .C(n65714), .D(
        \GFill[23][0] ), .S0(n65811), .S1(n65923), .Q(n14872) );
  IMUX40 U30572 ( .A(n65696), .B(n65697), .C(\GFill[38][0] ), .D(n65699), .S0(
        n65820), .S1(n65914), .Q(n25747) );
  IMUX40 U30568 ( .A(n65680), .B(n65681), .C(\GFill[54][0] ), .D(n65683), .S0(
        n65824), .S1(n65913), .Q(n25742) );
  IMUX40 U30580 ( .A(n65728), .B(\GFill[5][0] ), .C(n65730), .D(n65731), .S0(
        n65791), .S1(N1172), .Q(n25757) );
  IMUX40 U30576 ( .A(n65712), .B(n65713), .C(\GFill[22][0] ), .D(n65715), .S0(
        n65808), .S1(N1172), .Q(n25752) );
  IMUX40 U29900 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65883), .S1(n65752), .Q(n25107) );
  IMUX40 U29896 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65908), .S1(n65752), .Q(n25102) );
  IMUX40 U29908 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65868), .S1(n65753), .Q(n25117) );
  IMUX40 U29904 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65843), .S1(n65752), .Q(n25112) );
  IMUX40 U31244 ( .A(n65696), .B(n65697), .C(\GFill[38][0] ), .D(n65699), .S0(
        n65885), .S1(n65769), .Q(n26387) );
  IMUX40 U31240 ( .A(n65680), .B(n65681), .C(\GFill[54][0] ), .D(n65683), .S0(
        n65903), .S1(n65759), .Q(n26382) );
  IMUX40 U31252 ( .A(n65728), .B(\GFill[5][0] ), .C(n65730), .D(\GFill[7][0] ), 
        .S0(n65901), .S1(n65779), .Q(n26397) );
  IMUX40 U31248 ( .A(n65712), .B(n65713), .C(\GFill[22][0] ), .D(n65715), .S0(
        n65892), .S1(n65764), .Q(n26392) );
  IMUX40 U32588 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65790), .S1(n65537), .Q(n27667) );
  IMUX40 U32584 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65795), .S1(n65912), .Q(n27662) );
  IMUX40 U32596 ( .A(n65728), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(n65731), 
        .S0(n65805), .S1(N1130), .Q(n27677) );
  IMUX40 U32592 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65797), .S1(n65538), .Q(n27672) );
  IMUX40 U31916 ( .A(n65696), .B(n65697), .C(\GFill[38][0] ), .D(
        \GFill[39][0] ), .S0(n65864), .S1(n65777), .Q(n27027) );
  IMUX40 U31912 ( .A(n65680), .B(n65681), .C(\GFill[54][0] ), .D(
        \GFill[55][0] ), .S0(n65846), .S1(n65780), .Q(n27022) );
  IMUX40 U31924 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(n65730), .D(
        \GFill[7][0] ), .S0(n65884), .S1(n65771), .Q(n27037) );
  IMUX40 U31920 ( .A(n65712), .B(n65713), .C(\GFill[22][0] ), .D(
        \GFill[23][0] ), .S0(n65839), .S1(n65776), .Q(n27032) );
  IMUX40 U33260 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(n65699), .S0(n65866), .S1(n65744), .Q(n28307) );
  IMUX40 U33256 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(n65683), .S0(n65887), .S1(n65746), .Q(n28302) );
  IMUX40 U33268 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        n65731), .S0(n65842), .S1(n65744), .Q(n28317) );
  IMUX40 U33264 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(n65715), .S0(n65846), .S1(n65744), .Q(n28312) );
  IMUX40 U21836 ( .A(\GFill[36][0] ), .B(n65697), .C(n65698), .D(
        \GFill[39][0] ), .S0(n65847), .S1(n65773), .Q(n17427) );
  IMUX40 U21832 ( .A(\GFill[52][0] ), .B(n65681), .C(n65682), .D(
        \GFill[55][0] ), .S0(n65849), .S1(n65777), .Q(n17422) );
  IMUX40 U21844 ( .A(\GFill[4][0] ), .B(n65729), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65844), .S1(n65770), .Q(n17437) );
  IMUX40 U21840 ( .A(\GFill[20][0] ), .B(n65713), .C(n65714), .D(
        \GFill[23][0] ), .S0(n65846), .S1(n65776), .Q(n17432) );
  IMUX40 U23180 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65881), .S1(n65755), .Q(n18707) );
  IMUX40 U23176 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65836), .S1(n65754), .Q(n18702) );
  IMUX40 U23188 ( .A(n65728), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65906), .S1(N1208), .Q(n18717) );
  IMUX40 U23184 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65881), .S1(n65747), .Q(n18712) );
  IMUX40 U22508 ( .A(\GFill[36][0] ), .B(n65697), .C(n65698), .D(
        \GFill[39][0] ), .S0(n65793), .S1(N1172), .Q(n18067) );
  IMUX40 U22504 ( .A(\GFill[52][0] ), .B(n65681), .C(n65682), .D(
        \GFill[55][0] ), .S0(n65811), .S1(N1172), .Q(n18062) );
  IMUX40 U22516 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65785), .S1(N1172), .Q(n18077) );
  IMUX40 U22512 ( .A(\GFill[20][0] ), .B(n65713), .C(n65714), .D(
        \GFill[23][0] ), .S0(n65811), .S1(N1112), .Q(n18072) );
  IMUX40 U34604 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65805), 
        .S1(n65922), .Q(n29587) );
  IMUX40 U34600 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65800), 
        .S1(n65923), .Q(n29582) );
  IMUX40 U34612 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65809), 
        .S1(n65912), .Q(n29597) );
  IMUX40 U34608 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65808), 
        .S1(n65923), .Q(n29592) );
  IMUX40 U33932 ( .A(\GFill[36][0] ), .B(n65697), .C(n65698), .D(n65699), .S0(
        n65833), .S1(n65761), .Q(n28947) );
  IMUX40 U33928 ( .A(\GFill[52][0] ), .B(n65681), .C(n65682), .D(n65683), .S0(
        n65836), .S1(n65761), .Q(n28942) );
  IMUX40 U33940 ( .A(\GFill[4][0] ), .B(n65729), .C(n65730), .D(n65731), .S0(
        n65886), .S1(n65774), .Q(n28957) );
  IMUX40 U33936 ( .A(\GFill[20][0] ), .B(n65713), .C(n65714), .D(n65715), .S0(
        n65849), .S1(n65760), .Q(n28952) );
  IMUX40 U35276 ( .A(n65696), .B(n65697), .C(n65698), .D(n65699), .S0(n65867), 
        .S1(n65754), .Q(n30227) );
  IMUX40 U35272 ( .A(n65680), .B(n65681), .C(n65682), .D(n65683), .S0(n65881), 
        .S1(n65754), .Q(n30222) );
  IMUX40 U35284 ( .A(n65728), .B(n65729), .C(n65730), .D(n65731), .S0(n65875), 
        .S1(n65755), .Q(n30237) );
  IMUX40 U35280 ( .A(n65712), .B(n65713), .C(n65714), .D(n65715), .S0(n65842), 
        .S1(n65754), .Q(n30232) );
  IMUX40 U54764 ( .A(\OFill[36][0] ), .B(n65633), .C(n65634), .D(
        \OFill[39][0] ), .S0(n65791), .S1(N1112), .Q(n48787) );
  IMUX40 U54760 ( .A(\OFill[52][0] ), .B(n65617), .C(n65618), .D(
        \OFill[55][0] ), .S0(n65821), .S1(n65921), .Q(n48782) );
  IMUX40 U54772 ( .A(\OFill[4][0] ), .B(n65665), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65813), .S1(n65921), .Q(n48797) );
  IMUX40 U54768 ( .A(\OFill[20][0] ), .B(n65649), .C(n65650), .D(n65651), .S0(
        n65821), .S1(N1112), .Q(n48792) );
  IMUX40 U54092 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65852), .S1(n65778), .Q(n48147) );
  IMUX40 U54088 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65850), .S1(n65766), .Q(n48142) );
  IMUX40 U54100 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65867), .S1(n65772), .Q(n48157) );
  IMUX40 U54096 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65853), .S1(n65768), .Q(n48152) );
  IMUX40 U55436 ( .A(\OFill[36][0] ), .B(n65633), .C(n65634), .D(
        \OFill[39][0] ), .S0(n65845), .S1(n65748), .Q(n49427) );
  IMUX40 U55432 ( .A(\OFill[52][0] ), .B(n65617), .C(n65618), .D(
        \OFill[55][0] ), .S0(n65844), .S1(N1208), .Q(n49422) );
  IMUX40 U55444 ( .A(\OFill[4][0] ), .B(n65665), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65850), .S1(n65749), .Q(n49437) );
  IMUX40 U55440 ( .A(\OFill[20][0] ), .B(n65649), .C(n65650), .D(n65651), .S0(
        n65853), .S1(n65749), .Q(n49432) );
  IMUX40 U66860 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65828), 
        .S1(N1082), .Q(n60307) );
  IMUX40 U66856 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65820), 
        .S1(N860), .Q(n60302) );
  IMUX40 U66868 ( .A(\OFill[4][0] ), .B(n65665), .C(n65666), .D(n65667), .S0(
        n65794), .S1(n65743), .Q(n60317) );
  IMUX40 U66864 ( .A(\OFill[20][0] ), .B(n65649), .C(n65650), .D(n65651), .S0(
        n65816), .S1(n65743), .Q(n60312) );
  IMUX40 U66188 ( .A(\OFill[36][0] ), .B(n65633), .C(n65634), .D(n65635), .S0(
        n65880), .S1(n65763), .Q(n59667) );
  IMUX40 U66184 ( .A(\OFill[52][0] ), .B(n65617), .C(n65618), .D(n65619), .S0(
        n65881), .S1(n65762), .Q(n59662) );
  IMUX40 U66196 ( .A(\OFill[4][0] ), .B(n65665), .C(n65666), .D(n65667), .S0(
        n65862), .S1(n65764), .Q(n59677) );
  IMUX40 U66192 ( .A(\OFill[20][0] ), .B(n65649), .C(n65650), .D(n65651), .S0(
        n65884), .S1(n65763), .Q(n59672) );
  IMUX40 U67532 ( .A(n65632), .B(n65633), .C(n65634), .D(n65635), .S0(n65841), 
        .S1(n65747), .Q(n60947) );
  IMUX40 U67528 ( .A(n65616), .B(n65617), .C(n65618), .D(n65619), .S0(n65906), 
        .S1(n65747), .Q(n60942) );
  IMUX40 U67540 ( .A(n65664), .B(n65665), .C(n65666), .D(n65667), .S0(n65892), 
        .S1(n65746), .Q(n60957) );
  IMUX40 U67536 ( .A(n65648), .B(n65649), .C(n65650), .D(n65651), .S0(N1207), 
        .S1(n65747), .Q(n60952) );
  IMUX40 U7724 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(n65698), .D(
        \GFill[39][0] ), .S0(n65788), .S1(n65535), .Q(n3987) );
  IMUX40 U7720 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(n65682), .D(
        \GFill[55][0] ), .S0(n65788), .S1(n65535), .Q(n3982) );
  IMUX40 U7732 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65786), .S1(n65535), .Q(n3997) );
  IMUX40 U7728 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(n65714), .D(
        \GFill[23][0] ), .S0(n65787), .S1(n65535), .Q(n3992) );
  IMUX40 U9068 ( .A(n65696), .B(\GFill[37][0] ), .C(\GFill[38][0] ), .D(
        \GFill[39][0] ), .S0(n65811), .S1(N704), .Q(n5267) );
  IMUX40 U9064 ( .A(n65680), .B(\GFill[53][0] ), .C(\GFill[54][0] ), .D(
        \GFill[55][0] ), .S0(n65787), .S1(N704), .Q(n5262) );
  IMUX40 U9076 ( .A(\GFill[4][0] ), .B(n65729), .C(n65730), .D(\GFill[7][0] ), 
        .S0(n65810), .S1(N704), .Q(n5277) );
  IMUX40 U9072 ( .A(n65712), .B(\GFill[21][0] ), .C(\GFill[22][0] ), .D(
        \GFill[23][0] ), .S0(n65811), .S1(N704), .Q(n5272) );
  IMUX40 U8396 ( .A(n65696), .B(\GFill[37][0] ), .C(n65698), .D(\GFill[39][0] ), .S0(n65809), .S1(n65536), .Q(n4627) );
  IMUX40 U8392 ( .A(n65680), .B(\GFill[53][0] ), .C(n65682), .D(\GFill[55][0] ), .S0(n65810), .S1(n65536), .Q(n4622) );
  IMUX40 U8404 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65789), .S1(n65536), .Q(n4637) );
  IMUX40 U8400 ( .A(n65712), .B(\GFill[21][0] ), .C(n65714), .D(\GFill[23][0] ), .S0(n65820), .S1(n65536), .Q(n4632) );
  IMUX40 U10412 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65819), .S1(N716), .Q(n6547) );
  IMUX40 U10408 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65819), .S1(N716), .Q(n6542) );
  IMUX40 U10420 ( .A(\GFill[4][0] ), .B(n65729), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65817), .S1(N716), .Q(n6557) );
  IMUX40 U10416 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65818), .S1(N716), .Q(n6552) );
  IMUX40 U9740 ( .A(n65696), .B(\GFill[37][0] ), .C(n65698), .D(\GFill[39][0] ), .S0(n65800), .S1(n65935), .Q(n5907) );
  IMUX40 U9736 ( .A(n65680), .B(\GFill[53][0] ), .C(n65682), .D(\GFill[55][0] ), .S0(n65799), .S1(n65935), .Q(n5902) );
  IMUX40 U9748 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(n65730), .D(
        \GFill[7][0] ), .S0(n65798), .S1(N998), .Q(n5917) );
  IMUX40 U9744 ( .A(n65712), .B(\GFill[21][0] ), .C(n65714), .D(\GFill[23][0] ), .S0(n65798), .S1(n65935), .Q(n5912) );
  IMUX40 U11084 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65830), .S1(N722), .Q(n7187) );
  IMUX40 U11080 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65830), .S1(N722), .Q(n7182) );
  IMUX40 U11088 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65831), .S1(N722), .Q(n7192) );
  IMUX40 U12428 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65804), .S1(N1022), .Q(n8467) );
  IMUX40 U12424 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65804), .S1(n65930), .Q(n8462) );
  IMUX40 U12436 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(n65730), .D(
        \GFill[7][0] ), .S0(n65803), .S1(n65930), .Q(n8477) );
  IMUX40 U12432 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65802), .S1(n65932), .Q(n8472) );
  IMUX40 U11756 ( .A(n65696), .B(\GFill[37][0] ), .C(\GFill[38][0] ), .D(
        \GFill[39][0] ), .S0(n65808), .S1(n65933), .Q(n7827) );
  IMUX40 U11752 ( .A(n65680), .B(\GFill[53][0] ), .C(\GFill[54][0] ), .D(
        \GFill[55][0] ), .S0(n65828), .S1(n65930), .Q(n7822) );
  IMUX40 U11764 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65796), .S1(n65933), .Q(n7837) );
  IMUX40 U11760 ( .A(n65712), .B(\GFill[21][0] ), .C(\GFill[22][0] ), .D(
        \GFill[23][0] ), .S0(n65794), .S1(n65930), .Q(n7832) );
  IMUX40 U13100 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(n65699), .S0(n65823), .S1(N740), .Q(n9107) );
  IMUX40 U13096 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(n65683), .S0(n65823), .S1(N740), .Q(n9102) );
  IMUX40 U13108 ( .A(n65728), .B(\GFill[5][0] ), .C(n65730), .D(\GFill[7][0] ), 
        .S0(n65825), .S1(N740), .Q(n9117) );
  IMUX40 U13104 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(n65715), .S0(n65824), .S1(N740), .Q(n9112) );
  IMUX40 U13772 ( .A(n65696), .B(\GFill[37][0] ), .C(\GFill[38][0] ), .D(
        \GFill[39][0] ), .S0(n65792), .S1(n65929), .Q(n9747) );
  IMUX40 U13768 ( .A(n65680), .B(\GFill[53][0] ), .C(\GFill[54][0] ), .D(
        \GFill[55][0] ), .S0(n65791), .S1(n65929), .Q(n9742) );
  IMUX40 U13780 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        n65731), .S0(n65790), .S1(N1034), .Q(n9757) );
  IMUX40 U13776 ( .A(n65712), .B(\GFill[21][0] ), .C(\GFill[22][0] ), .D(
        \GFill[23][0] ), .S0(n65789), .S1(n65929), .Q(n9752) );
  IMUX40 U15116 ( .A(\GFill[36][0] ), .B(n65697), .C(\GFill[38][0] ), .D(
        n65699), .S0(n65796), .S1(n65925), .Q(n11027) );
  IMUX40 U15112 ( .A(\GFill[52][0] ), .B(n65681), .C(\GFill[54][0] ), .D(
        n65683), .S0(n65796), .S1(N1010), .Q(n11022) );
  IMUX40 U15124 ( .A(n65728), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65794), .S1(N1010), .Q(n11037) );
  IMUX40 U15120 ( .A(\GFill[20][0] ), .B(n65713), .C(\GFill[22][0] ), .D(
        n65715), .S0(n65794), .S1(N1046), .Q(n11032) );
  IMUX40 U14444 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65823), .S1(n65927), .Q(n10387) );
  IMUX40 U14440 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65807), .S1(n65927), .Q(n10382) );
  IMUX40 U14452 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        n65731), .S0(n65783), .S1(N1040), .Q(n10397) );
  IMUX40 U14448 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65826), .S1(n65927), .Q(n10392) );
  IMUX40 U28556 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(n65699), .S0(n65880), .S1(n65751), .Q(n23827) );
  IMUX40 U28552 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(n65683), .S0(n65906), .S1(n65751), .Q(n23822) );
  IMUX40 U28564 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        n65731), .S0(n65883), .S1(n65751), .Q(n23837) );
  IMUX40 U28560 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(n65715), .S0(n65871), .S1(n65751), .Q(n23832) );
  IMUX40 U27884 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65874), .S1(n65772), .Q(n23187) );
  IMUX40 U27880 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65896), .S1(n65759), .Q(n23182) );
  IMUX40 U27892 ( .A(n65728), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65882), .S1(n65769), .Q(n23197) );
  IMUX40 U27888 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65876), .S1(n65776), .Q(n23192) );
  IMUX40 U29228 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(n65699), .S0(n65792), .S1(n65913), .Q(n24467) );
  IMUX40 U29224 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(n65683), .S0(n65808), .S1(N1184), .Q(n24462) );
  IMUX40 U29236 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65798), .S1(n65913), .Q(n24477) );
  IMUX40 U29232 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(n65715), .S0(n65799), .S1(N1184), .Q(n24472) );
  IMUX40 U26540 ( .A(n65696), .B(\GFill[37][0] ), .C(\GFill[38][0] ), .D(
        \GFill[39][0] ), .S0(n65788), .S1(n65534), .Q(n21907) );
  IMUX40 U26536 ( .A(n65680), .B(\GFill[53][0] ), .C(\GFill[54][0] ), .D(
        \GFill[55][0] ), .S0(n65783), .S1(n65534), .Q(n21902) );
  IMUX40 U26548 ( .A(n65728), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(n65731), 
        .S0(n65797), .S1(n65534), .Q(n21917) );
  IMUX40 U26544 ( .A(n65712), .B(\GFill[21][0] ), .C(\GFill[22][0] ), .D(
        \GFill[23][0] ), .S0(n65796), .S1(n65534), .Q(n21912) );
  IMUX40 U25868 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(n65698), .D(
        \GFill[39][0] ), .S0(n65886), .S1(n65759), .Q(n21267) );
  IMUX40 U25864 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(n65682), .D(
        \GFill[55][0] ), .S0(n65885), .S1(n65781), .Q(n21262) );
  IMUX40 U25876 ( .A(\GFill[4][0] ), .B(n65729), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65880), .S1(n65762), .Q(n21277) );
  IMUX40 U25872 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(n65714), .D(
        \GFill[23][0] ), .S0(n65907), .S1(n65777), .Q(n21272) );
  IMUX40 U27212 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65841), .S1(n65746), .Q(n22547) );
  IMUX40 U27208 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65870), .S1(n65745), .Q(n22542) );
  IMUX40 U27220 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65838), .S1(n65746), .Q(n22557) );
  IMUX40 U27216 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65905), .S1(n65746), .Q(n22552) );
  IMUX40 U24524 ( .A(n65696), .B(\GFill[37][0] ), .C(\GFill[38][0] ), .D(
        \GFill[39][0] ), .S0(n65799), .S1(N842), .Q(n19987) );
  IMUX40 U24520 ( .A(n65680), .B(\GFill[53][0] ), .C(\GFill[54][0] ), .D(
        \GFill[55][0] ), .S0(n65829), .S1(N842), .Q(n19982) );
  IMUX40 U24532 ( .A(\GFill[4][0] ), .B(n65729), .C(n65730), .D(\GFill[7][0] ), 
        .S0(n65824), .S1(N842), .Q(n19997) );
  IMUX40 U24528 ( .A(n65712), .B(\GFill[21][0] ), .C(\GFill[22][0] ), .D(
        \GFill[23][0] ), .S0(n65784), .S1(N842), .Q(n19992) );
  IMUX40 U23852 ( .A(\GFill[36][0] ), .B(\GFill[37][0] ), .C(\GFill[38][0] ), 
        .D(\GFill[39][0] ), .S0(n65899), .S1(n65764), .Q(n19347) );
  IMUX40 U23848 ( .A(\GFill[52][0] ), .B(\GFill[53][0] ), .C(\GFill[54][0] ), 
        .D(\GFill[55][0] ), .S0(n65843), .S1(n65776), .Q(n19342) );
  IMUX40 U23860 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(\GFill[6][0] ), .D(
        \GFill[7][0] ), .S0(n65901), .S1(n65773), .Q(n19357) );
  IMUX40 U23856 ( .A(\GFill[20][0] ), .B(\GFill[21][0] ), .C(\GFill[22][0] ), 
        .D(\GFill[23][0] ), .S0(n65836), .S1(n65766), .Q(n19352) );
  IMUX40 U25196 ( .A(n65696), .B(\GFill[37][0] ), .C(\GFill[38][0] ), .D(
        \GFill[39][0] ), .S0(n65854), .S1(n65744), .Q(n20627) );
  IMUX40 U25192 ( .A(n65680), .B(\GFill[53][0] ), .C(\GFill[54][0] ), .D(
        \GFill[55][0] ), .S0(n65855), .S1(n65746), .Q(n20622) );
  IMUX40 U25204 ( .A(\GFill[4][0] ), .B(\GFill[5][0] ), .C(n65730), .D(
        \GFill[7][0] ), .S0(n65893), .S1(n65754), .Q(n20637) );
  IMUX40 U25200 ( .A(n65712), .B(\GFill[21][0] ), .C(\GFill[22][0] ), .D(
        \GFill[23][0] ), .S0(n65856), .S1(n65753), .Q(n20632) );
  IMUX40 U40652 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(n65634), .D(
        \OFill[39][0] ), .S0(n65814), .S1(n65924), .Q(n35347) );
  IMUX40 U40648 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(n65618), .D(
        \OFill[55][0] ), .S0(n65815), .S1(N980), .Q(n35342) );
  IMUX40 U40660 ( .A(\OFill[4][0] ), .B(n65665), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65813), .S1(N1010), .Q(n35357) );
  IMUX40 U40656 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(n65650), .D(
        n65651), .S0(n65813), .S1(n65925), .Q(n35352) );
  IMUX40 U39980 ( .A(n65632), .B(\OFill[37][0] ), .C(\OFill[38][0] ), .D(
        \OFill[39][0] ), .S0(n65812), .S1(N1046), .Q(n34707) );
  IMUX40 U39976 ( .A(n65616), .B(\OFill[53][0] ), .C(\OFill[54][0] ), .D(
        \OFill[55][0] ), .S0(n65812), .S1(N1046), .Q(n34702) );
  IMUX40 U39988 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65804), .S1(N1046), .Q(n34717) );
  IMUX40 U39984 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65821), .S1(N1046), .Q(n34712) );
  IMUX40 U41324 ( .A(n65632), .B(\OFill[37][0] ), .C(n65634), .D(
        \OFill[39][0] ), .S0(n65816), .S1(N1004), .Q(n35987) );
  IMUX40 U41320 ( .A(n65616), .B(\OFill[53][0] ), .C(n65618), .D(
        \OFill[55][0] ), .S0(n65817), .S1(N1004), .Q(n35982) );
  IMUX40 U41332 ( .A(n65664), .B(n65665), .C(\OFill[6][0] ), .D(\OFill[7][0] ), 
        .S0(n65815), .S1(N1004), .Q(n35997) );
  IMUX40 U41328 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(n65650), .D(
        n65651), .S0(n65816), .S1(N1004), .Q(n35992) );
  IMUX40 U42668 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65828), .S1(N1034), .Q(n37267) );
  IMUX40 U42664 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65828), .S1(N1034), .Q(n37262) );
  IMUX40 U42676 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65830), .S1(N1034), .Q(n37277) );
  IMUX40 U42672 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65829), .S1(N1034), .Q(n37272) );
  IMUX40 U41996 ( .A(n65632), .B(\OFill[37][0] ), .C(n65634), .D(
        \OFill[39][0] ), .S0(n65801), .S1(n65934), .Q(n36627) );
  IMUX40 U41992 ( .A(n65616), .B(\OFill[53][0] ), .C(n65618), .D(
        \OFill[55][0] ), .S0(n65798), .S1(n65935), .Q(n36622) );
  IMUX40 U42004 ( .A(n65664), .B(n65665), .C(\OFill[6][0] ), .D(\OFill[7][0] ), 
        .S0(n65800), .S1(n65934), .Q(n36637) );
  IMUX40 U42000 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(n65650), .D(
        n65651), .S0(n65801), .S1(n65934), .Q(n36632) );
  IMUX40 U43340 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65826), .S1(n65925), .Q(n37907) );
  IMUX40 U43336 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65825), .S1(n65924), .Q(n37902) );
  IMUX40 U43348 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65827), .S1(N1010), .Q(n37917) );
  IMUX40 U43344 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65826), .S1(N980), .Q(n37912) );
  IMUX40 U44684 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65806), .S1(n65932), .Q(n39187) );
  IMUX40 U44680 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65803), .S1(n65930), .Q(n39182) );
  IMUX40 U44692 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65805), .S1(n65932), .Q(n39197) );
  IMUX40 U44688 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65805), .S1(n65931), .Q(n39192) );
  IMUX40 U44012 ( .A(n65632), .B(\OFill[37][0] ), .C(\OFill[38][0] ), .D(
        \OFill[39][0] ), .S0(n65814), .S1(n65932), .Q(n38547) );
  IMUX40 U44008 ( .A(n65616), .B(\OFill[53][0] ), .C(\OFill[54][0] ), .D(
        \OFill[55][0] ), .S0(n65820), .S1(n65932), .Q(n38542) );
  IMUX40 U44020 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65809), .S1(n65931), .Q(n38557) );
  IMUX40 U44016 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65815), .S1(n65931), .Q(n38552) );
  IMUX40 U45356 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(n65635), .S0(n65826), .S1(N1040), .Q(n39827) );
  IMUX40 U45352 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(n65619), .S0(n65821), .S1(N1040), .Q(n39822) );
  IMUX40 U45364 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        n65667), .S0(n65822), .S1(N1040), .Q(n39837) );
  IMUX40 U45360 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65822), .S1(N1040), .Q(n39832) );
  IMUX40 U46700 ( .A(n65632), .B(\OFill[37][0] ), .C(\OFill[38][0] ), .D(
        \OFill[39][0] ), .S0(n65782), .S1(n65926), .Q(n41107) );
  IMUX40 U46696 ( .A(n65616), .B(\OFill[53][0] ), .C(\OFill[54][0] ), .D(
        \OFill[55][0] ), .S0(n65819), .S1(n65927), .Q(n41102) );
  IMUX40 U46708 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65807), .S1(n65926), .Q(n41117) );
  IMUX40 U46704 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65794), .S1(n65926), .Q(n41112) );
  IMUX40 U46028 ( .A(\OFill[36][0] ), .B(n65633), .C(\OFill[38][0] ), .D(
        n65635), .S0(n65793), .S1(n65928), .Q(n40467) );
  IMUX40 U46024 ( .A(\OFill[52][0] ), .B(n65617), .C(\OFill[54][0] ), .D(
        n65619), .S0(n65790), .S1(n65929), .Q(n40462) );
  IMUX40 U46036 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(n65666), .D(n65667), 
        .S0(n65792), .S1(n65928), .Q(n40477) );
  IMUX40 U46032 ( .A(\OFill[20][0] ), .B(n65649), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65793), .S1(n65928), .Q(n40472) );
  IMUX40 U47372 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65812), .S1(n65925), .Q(n41747) );
  IMUX40 U47368 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65795), .S1(n65925), .Q(n41742) );
  IMUX40 U47380 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65797), .S1(n65924), .Q(n41757) );
  IMUX40 U47376 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65797), .S1(n65924), .Q(n41752) );
  IMUX40 U60812 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(n65635), .S0(n65907), .S1(n65750), .Q(n54547) );
  IMUX40 U60808 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(n65619), .S0(n65859), .S1(n65750), .Q(n54542) );
  IMUX40 U60820 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(n65666), .D(n65667), 
        .S0(n65848), .S1(n65749), .Q(n54557) );
  IMUX40 U60816 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65899), .S1(n65750), .Q(n54552) );
  IMUX40 U60140 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65856), .S1(n65770), .Q(n53907) );
  IMUX40 U60136 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65834), .S1(n65777), .Q(n53902) );
  IMUX40 U60148 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65883), .S1(n65781), .Q(n53917) );
  IMUX40 U60144 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65909), .S1(n65771), .Q(n53912) );
  IMUX40 U61484 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(n65635), .S0(n65824), .S1(N1172), .Q(n55187) );
  IMUX40 U61480 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(n65619), .S0(n65823), .S1(n65914), .Q(n55182) );
  IMUX40 U61492 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(n65666), .D(n65667), 
        .S0(n65787), .S1(n65914), .Q(n55197) );
  IMUX40 U61488 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(n65651), .S0(n65788), .S1(N1184), .Q(n55192) );
  IMUX40 U58796 ( .A(n65632), .B(\OFill[37][0] ), .C(\OFill[38][0] ), .D(
        \OFill[39][0] ), .S0(n65796), .S1(n65537), .Q(n52627) );
  IMUX40 U58792 ( .A(n65616), .B(\OFill[53][0] ), .C(\OFill[54][0] ), .D(
        \OFill[55][0] ), .S0(n65794), .S1(n65911), .Q(n52622) );
  IMUX40 U58804 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65820), .S1(n65537), .Q(n52637) );
  IMUX40 U58800 ( .A(n65648), .B(\OFill[21][0] ), .C(\OFill[22][0] ), .D(
        \OFill[23][0] ), .S0(n65830), .S1(n65537), .Q(n52632) );
  IMUX40 U58124 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(n65634), .D(
        \OFill[39][0] ), .S0(n65904), .S1(n65773), .Q(n51987) );
  IMUX40 U58120 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(n65618), .D(
        \OFill[55][0] ), .S0(n65872), .S1(n65776), .Q(n51982) );
  IMUX40 U58132 ( .A(\OFill[4][0] ), .B(n65665), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65875), .S1(n65778), .Q(n51997) );
  IMUX40 U58128 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(n65650), .D(
        n65651), .S0(n65887), .S1(n65781), .Q(n51992) );
  IMUX40 U59468 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65844), .S1(n65745), .Q(n53267) );
  IMUX40 U59464 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65893), .S1(n65745), .Q(n53262) );
  IMUX40 U59476 ( .A(n65664), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65883), .S1(n65744), .Q(n53277) );
  IMUX40 U59472 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65875), .S1(n65744), .Q(n53272) );
  IMUX40 U56780 ( .A(n65632), .B(\OFill[37][0] ), .C(\OFill[38][0] ), .D(
        \OFill[39][0] ), .S0(n65784), .S1(n65912), .Q(n50707) );
  IMUX40 U56776 ( .A(n65616), .B(\OFill[53][0] ), .C(\OFill[54][0] ), .D(
        \OFill[55][0] ), .S0(n65785), .S1(n65923), .Q(n50702) );
  IMUX40 U56788 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65783), .S1(n65538), .Q(n50717) );
  IMUX40 U56784 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65784), .S1(n65538), .Q(n50712) );
  IMUX40 U56108 ( .A(\OFill[36][0] ), .B(\OFill[37][0] ), .C(\OFill[38][0] ), 
        .D(\OFill[39][0] ), .S0(n65878), .S1(n65771), .Q(n50067) );
  IMUX40 U56104 ( .A(\OFill[52][0] ), .B(\OFill[53][0] ), .C(\OFill[54][0] ), 
        .D(\OFill[55][0] ), .S0(n65834), .S1(n65775), .Q(n50062) );
  IMUX40 U56116 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65902), .S1(n65774), .Q(n50077) );
  IMUX40 U56112 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65890), .S1(n65771), .Q(n50072) );
  IMUX40 U57452 ( .A(n65632), .B(\OFill[37][0] ), .C(\OFill[38][0] ), .D(
        \OFill[39][0] ), .S0(n65884), .S1(n65748), .Q(n51347) );
  IMUX40 U57448 ( .A(n65616), .B(\OFill[53][0] ), .C(\OFill[54][0] ), .D(
        \OFill[55][0] ), .S0(N1207), .S1(n65748), .Q(n51342) );
  IMUX40 U57460 ( .A(\OFill[4][0] ), .B(\OFill[5][0] ), .C(\OFill[6][0] ), .D(
        \OFill[7][0] ), .S0(n65870), .S1(n65748), .Q(n51357) );
  IMUX40 U57456 ( .A(\OFill[20][0] ), .B(\OFill[21][0] ), .C(\OFill[22][0] ), 
        .D(\OFill[23][0] ), .S0(n65834), .S1(n65748), .Q(n51352) );
  IMUX40 U62833 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(n65646), .D(
        n65647), .S0(n65829), .S1(n65913), .Q(n56470) );
  IMUX40 U62830 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(n65659), .S0(n65806), .S1(N1184), .Q(n56473) );
  IMUX40 U62831 ( .A(\OFill[24][0] ), .B(n65653), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65827), .S1(N1172), .Q(n56471) );
  IMUX40 U62664 ( .A(n56470), .B(n56471), .C(n56472), .D(n56473), .S0(N1186), 
        .S1(N1185), .Q(n56469) );
  IMUX40 U30577 ( .A(n65708), .B(n65709), .C(\GFill[18][0] ), .D(n65711), .S0(
        n65801), .S1(n65913), .Q(n25750) );
  IMUX40 U30574 ( .A(n65720), .B(n65721), .C(\GFill[30][0] ), .D(n65723), .S0(
        n65791), .S1(n65913), .Q(n25753) );
  IMUX40 U30575 ( .A(n65716), .B(n65717), .C(\GFill[26][0] ), .D(n65719), .S0(
        n65787), .S1(N1184), .Q(n25751) );
  IMUX40 U30408 ( .A(n25750), .B(n25751), .C(n25752), .D(n25753), .S0(N1186), 
        .S1(N1185), .Q(n25749) );
  IMUX40 U22513 ( .A(n65708), .B(\GFill[17][0] ), .C(\GFill[18][0] ), .D(
        \GFill[19][0] ), .S0(n65785), .S1(N1112), .Q(n18070) );
  IMUX40 U22510 ( .A(n65720), .B(\GFill[29][0] ), .C(\GFill[30][0] ), .D(
        \GFill[31][0] ), .S0(n65807), .S1(n65921), .Q(n18073) );
  IMUX40 U22511 ( .A(n65716), .B(\GFill[25][0] ), .C(\GFill[26][0] ), .D(
        \GFill[27][0] ), .S0(n65784), .S1(n65913), .Q(n18071) );
  IMUX40 U22344 ( .A(n18070), .B(n18071), .C(n18072), .D(n18073), .S0(N1114), 
        .S1(N1113), .Q(n18069) );
  IMUX40 U54773 ( .A(n65660), .B(n65661), .C(\OFill[2][0] ), .D(\OFill[3][0] ), 
        .S0(n65783), .S1(n65921), .Q(n48795) );
  IMUX40 U54770 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65802), .S1(n65921), .Q(n48798) );
  IMUX40 U54771 ( .A(\OFill[8][0] ), .B(n65669), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65812), .S1(N1112), .Q(n48796) );
  IMUX40 U54601 ( .A(n48795), .B(n48796), .C(n48797), .D(n48798), .S0(N1114), 
        .S1(N1113), .Q(n48794) );
  IMUX40 U54769 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65801), .S1(n65921), .Q(n48790) );
  IMUX40 U54766 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65799), .S1(N1112), .Q(n48793) );
  IMUX40 U54767 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65798), .S1(n65921), .Q(n48791) );
  IMUX40 U54600 ( .A(n48790), .B(n48791), .C(n48792), .D(n48793), .S0(N1114), 
        .S1(N1113), .Q(n48789) );
  IMUX40 U7733 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65786), .S1(n65535), .Q(n3995) );
  IMUX40 U7730 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65787), .S1(n65535), .Q(n3998) );
  IMUX40 U7731 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(
        \GFill[11][0] ), .S0(n65787), .S1(n65535), .Q(n3996) );
  IMUX40 U7561 ( .A(n3995), .B(n3996), .C(n3997), .D(n3998), .S0(N694), .S1(
        N693), .Q(n3994) );
  IMUX40 U7729 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(n65710), .D(
        \GFill[19][0] ), .S0(n65787), .S1(n65535), .Q(n3990) );
  IMUX40 U7726 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(n65722), .D(
        \GFill[31][0] ), .S0(n65787), .S1(n65535), .Q(n3993) );
  IMUX40 U7727 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(n65718), .D(
        \GFill[27][0] ), .S0(n65787), .S1(n65535), .Q(n3991) );
  IMUX40 U7560 ( .A(n3990), .B(n3991), .C(n3992), .D(n3993), .S0(N694), .S1(
        N693), .Q(n3989) );
  IMUX40 U8401 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65789), .S1(n65536), .Q(n4630) );
  IMUX40 U8398 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65809), .S1(n65536), .Q(n4633) );
  IMUX40 U8399 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65809), .S1(n65536), .Q(n4631) );
  IMUX40 U8232 ( .A(n4630), .B(n4631), .C(n4632), .D(n4633), .S0(N700), .S1(
        N699), .Q(n4629) );
  IMUX40 U29233 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65806), .S1(n65914), .Q(n24470) );
  IMUX40 U29230 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65793), .S1(n65914), .Q(n24473) );
  IMUX40 U29231 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65801), .S1(N1172), .Q(n24471) );
  IMUX40 U29064 ( .A(n24470), .B(n24471), .C(n24472), .D(n24473), .S0(N1174), 
        .S1(N1173), .Q(n24469) );
  IMUX40 U24529 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(n65711), .S0(n65789), .S1(N842), .Q(n19990) );
  IMUX40 U24526 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(n65723), .S0(n65831), .S1(N842), .Q(n19993) );
  IMUX40 U24527 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(n65719), .S0(n65811), .S1(N842), .Q(n19991) );
  IMUX40 U24360 ( .A(n19990), .B(n19991), .C(n19992), .D(n19993), .S0(N844), 
        .S1(N843), .Q(n19989) );
  IMUX40 U70897 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65784), 
        .S1(N1256), .Q(n64150) );
  IMUX40 U70894 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65782), 
        .S1(N1256), .Q(n64153) );
  IMUX40 U70895 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65801), 
        .S1(N1256), .Q(n64151) );
  IMUX40 U70728 ( .A(n64150), .B(n64151), .C(n64152), .D(n64153), .S0(N1258), 
        .S1(N1257), .Q(n64149) );
  IMUX40 U61489 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65801), .S1(N1172), .Q(n55190) );
  IMUX40 U61486 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65815), .S1(N1112), .Q(n55193) );
  IMUX40 U61487 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65807), .S1(n65914), .Q(n55191) );
  IMUX40 U61320 ( .A(n55190), .B(n55191), .C(n55192), .D(n55193), .S0(N1174), 
        .S1(N1173), .Q(n55189) );
  IMUX40 U38641 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65788), 
        .S1(N968), .Q(n33430) );
  IMUX40 U38638 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65783), 
        .S1(N968), .Q(n33433) );
  IMUX40 U38639 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65793), 
        .S1(N968), .Q(n33431) );
  IMUX40 U38472 ( .A(n33430), .B(n33431), .C(n33432), .D(n33433), .S0(N970), 
        .S1(N969), .Q(n33429) );
  IMUX40 U37301 ( .A(n65724), .B(n65725), .C(n65726), .D(n65727), .S0(n65786), 
        .S1(N956), .Q(n32155) );
  IMUX40 U37298 ( .A(n65736), .B(n65737), .C(n65738), .D(n65739), .S0(n65793), 
        .S1(N956), .Q(n32158) );
  IMUX40 U37299 ( .A(n65732), .B(n65733), .C(n65734), .D(n65735), .S0(n65792), 
        .S1(N956), .Q(n32156) );
  IMUX40 U37129 ( .A(n32155), .B(n32156), .C(n32157), .D(n32158), .S0(N958), 
        .S1(N957), .Q(n32154) );
  IMUX40 U69557 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65788), 
        .S1(N1244), .Q(n62875) );
  IMUX40 U69555 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65831), 
        .S1(N1244), .Q(n62876) );
  IMUX40 U69554 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65820), 
        .S1(N1244), .Q(n62878) );
  IMUX40 U69385 ( .A(n62875), .B(n62876), .C(n62877), .D(n62878), .S0(N1246), 
        .S1(N1245), .Q(n62874) );
  IMUX40 U13101 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65824), .S1(N740), .Q(n9105) );
  IMUX40 U13098 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65823), .S1(N740), .Q(n9108) );
  IMUX40 U13099 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65823), .S1(N740), .Q(n9106) );
  IMUX40 U12935 ( .A(n9105), .B(n9106), .C(n9107), .D(n9108), .S0(N742), .S1(
        N741), .Q(n9104) );
  IMUX40 U13097 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65823), .S1(N740), .Q(n9100) );
  IMUX40 U13094 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65823), .S1(N740), .Q(n9103) );
  IMUX40 U13095 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65823), .S1(N740), .Q(n9101) );
  IMUX40 U12934 ( .A(n9100), .B(n9101), .C(n9102), .D(n9103), .S0(N742), .S1(
        N741), .Q(n9099) );
  IMUX40 U40653 ( .A(n65628), .B(n65629), .C(\OFill[34][0] ), .D(n65631), .S0(
        n65814), .S1(N1010), .Q(n35345) );
  IMUX40 U40650 ( .A(n65640), .B(n65641), .C(\OFill[46][0] ), .D(n65643), .S0(
        n65814), .S1(N980), .Q(n35348) );
  IMUX40 U40651 ( .A(n65636), .B(n65637), .C(\OFill[42][0] ), .D(n65639), .S0(
        n65814), .S1(n65924), .Q(n35346) );
  IMUX40 U40487 ( .A(n35345), .B(n35346), .C(n35347), .D(n35348), .S0(N988), 
        .S1(N987), .Q(n35344) );
  IMUX40 U40649 ( .A(n65612), .B(n65613), .C(\OFill[50][0] ), .D(n65615), .S0(
        n65814), .S1(N980), .Q(n35340) );
  IMUX40 U40646 ( .A(n65624), .B(n65625), .C(\OFill[62][0] ), .D(n65627), .S0(
        n65815), .S1(N980), .Q(n35343) );
  IMUX40 U40647 ( .A(n65620), .B(n65621), .C(\OFill[58][0] ), .D(n65623), .S0(
        n65815), .S1(N980), .Q(n35341) );
  IMUX40 U40486 ( .A(n35340), .B(n35341), .C(n35342), .D(n35343), .S0(N988), 
        .S1(N987), .Q(n35339) );
  IMUX40 U39981 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65812), .S1(N1046), .Q(n34705) );
  IMUX40 U39978 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65812), .S1(N1046), .Q(n34708) );
  IMUX40 U39979 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65812), .S1(N1046), .Q(n34706) );
  IMUX40 U39815 ( .A(n34705), .B(n34706), .C(n34707), .D(n34708), .S0(N982), 
        .S1(N981), .Q(n34704) );
  IMUX40 U39977 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65812), .S1(N1046), .Q(n34700) );
  IMUX40 U39974 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65813), .S1(N1046), .Q(n34703) );
  IMUX40 U39975 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65812), .S1(N1046), .Q(n34701) );
  IMUX40 U39814 ( .A(n34700), .B(n34701), .C(n34702), .D(n34703), .S0(N982), 
        .S1(N981), .Q(n34699) );
  IMUX40 U26541 ( .A(\GFill[32][0] ), .B(n65693), .C(\GFill[34][0] ), .D(
        n65695), .S0(n65782), .S1(n65534), .Q(n21905) );
  IMUX40 U26538 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(n65706), .D(
        \GFill[47][0] ), .S0(n65789), .S1(n65534), .Q(n21908) );
  IMUX40 U26539 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(n65702), .D(
        \GFill[43][0] ), .S0(n65831), .S1(n65534), .Q(n21906) );
  IMUX40 U26375 ( .A(n21905), .B(n21906), .C(n21907), .D(n21908), .S0(N862), 
        .S1(N861), .Q(n21904) );
  IMUX40 U26537 ( .A(\GFill[48][0] ), .B(n65677), .C(\GFill[50][0] ), .D(
        n65679), .S0(n65783), .S1(n65534), .Q(n21900) );
  IMUX40 U26534 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(n65690), .D(
        \GFill[63][0] ), .S0(n65783), .S1(n65534), .Q(n21903) );
  IMUX40 U26535 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(n65686), .D(
        \GFill[59][0] ), .S0(n65783), .S1(n65534), .Q(n21901) );
  IMUX40 U26374 ( .A(n21900), .B(n21901), .C(n21902), .D(n21903), .S0(N862), 
        .S1(N861), .Q(n21899) );
  IMUX40 U58797 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65814), .S1(n65537), .Q(n52625) );
  IMUX40 U58794 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65793), .S1(n65922), .Q(n52628) );
  IMUX40 U58795 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65792), .S1(N1082), .Q(n52626) );
  IMUX40 U58631 ( .A(n52625), .B(n52626), .C(n52627), .D(n52628), .S0(N1150), 
        .S1(N1149), .Q(n52624) );
  IMUX40 U58793 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65827), .S1(N1082), .Q(n52620) );
  IMUX40 U58790 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65822), .S1(n65537), .Q(n52623) );
  IMUX40 U58791 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65815), .S1(n65538), .Q(n52621) );
  IMUX40 U58630 ( .A(n52620), .B(n52621), .C(n52622), .D(n52623), .S0(N1150), 
        .S1(N1149), .Q(n52619) );
  IMUX40 U56781 ( .A(n65628), .B(n65629), .C(n65630), .D(\OFill[35][0] ), .S0(
        n65784), .S1(N1082), .Q(n50705) );
  IMUX40 U56778 ( .A(n65640), .B(n65641), .C(n65642), .D(\OFill[47][0] ), .S0(
        n65785), .S1(n65537), .Q(n50708) );
  IMUX40 U56779 ( .A(n65636), .B(n65637), .C(n65638), .D(\OFill[43][0] ), .S0(
        n65785), .S1(N1082), .Q(n50706) );
  IMUX40 U56615 ( .A(n50705), .B(n50706), .C(n50707), .D(n50708), .S0(N1132), 
        .S1(N1131), .Q(n50704) );
  IMUX40 U56777 ( .A(n65612), .B(n65613), .C(n65614), .D(\OFill[51][0] ), .S0(
        n65785), .S1(n65911), .Q(n50700) );
  IMUX40 U56774 ( .A(n65624), .B(n65625), .C(n65626), .D(\OFill[63][0] ), .S0(
        n65785), .S1(n65912), .Q(n50703) );
  IMUX40 U56775 ( .A(n65620), .B(n65621), .C(n65622), .D(\OFill[59][0] ), .S0(
        n65785), .S1(n65743), .Q(n50701) );
  IMUX40 U56614 ( .A(n50700), .B(n50701), .C(n50702), .D(n50703), .S0(N1132), 
        .S1(N1131), .Q(n50699) );
  IMUX40 U39309 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(n65902), 
        .S1(n65768), .Q(n34065) );
  IMUX40 U39306 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65843), 
        .S1(n65768), .Q(n34068) );
  IMUX40 U39307 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65875), 
        .S1(n65768), .Q(n34066) );
  IMUX40 U39143 ( .A(n34065), .B(n34066), .C(n34067), .D(n34068), .S0(N976), 
        .S1(N975), .Q(n34064) );
  IMUX40 U39305 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65861), 
        .S1(n65767), .Q(n34060) );
  IMUX40 U39302 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(n65868), 
        .S1(n65767), .Q(n34063) );
  IMUX40 U39303 ( .A(n65684), .B(n65685), .C(n65686), .D(n65687), .S0(n65893), 
        .S1(n65767), .Q(n34061) );
  IMUX40 U39142 ( .A(n34060), .B(n34061), .C(n34062), .D(n34063), .S0(N976), 
        .S1(N975), .Q(n34059) );
  IMUX40 U36621 ( .A(n65692), .B(n65693), .C(n65694), .D(n65695), .S0(N1207), 
        .S1(n65755), .Q(n31505) );
  IMUX40 U36618 ( .A(n65704), .B(n65705), .C(n65706), .D(n65707), .S0(n65848), 
        .S1(n65756), .Q(n31508) );
  IMUX40 U36619 ( .A(n65700), .B(n65701), .C(n65702), .D(n65703), .S0(n65896), 
        .S1(n65755), .Q(n31506) );
  IMUX40 U36455 ( .A(n31505), .B(n31506), .C(n31507), .D(n31508), .S0(N952), 
        .S1(n65918), .Q(n31504) );
  IMUX40 U36617 ( .A(n65676), .B(n65677), .C(n65678), .D(n65679), .S0(n65847), 
        .S1(n65755), .Q(n31500) );
  IMUX40 U36614 ( .A(n65688), .B(n65689), .C(n65690), .D(n65691), .S0(n65853), 
        .S1(n65755), .Q(n31503) );
  IMUX40 U36615 ( .A(n65684), .B(n65685), .C(n65686), .D(n65687), .S0(n65910), 
        .S1(n65755), .Q(n31501) );
  IMUX40 U36454 ( .A(n31500), .B(n31501), .C(n31502), .D(n31503), .S0(N952), 
        .S1(n65917), .Q(n31499) );
  IMUX40 U68877 ( .A(n65628), .B(n65629), .C(n65630), .D(n65631), .S0(n65898), 
        .S1(n65749), .Q(n62225) );
  IMUX40 U68874 ( .A(n65640), .B(n65641), .C(n65642), .D(n65643), .S0(n65854), 
        .S1(n65756), .Q(n62228) );
  IMUX40 U68875 ( .A(n65636), .B(n65637), .C(n65638), .D(n65639), .S0(n65895), 
        .S1(n65756), .Q(n62226) );
  IMUX40 U68711 ( .A(n62225), .B(n62226), .C(n62227), .D(n62228), .S0(N1240), 
        .S1(n65918), .Q(n62224) );
  IMUX40 U68873 ( .A(n65612), .B(n65613), .C(n65614), .D(n65615), .S0(n65887), 
        .S1(n65756), .Q(n62220) );
  IMUX40 U68870 ( .A(n65624), .B(n65625), .C(n65626), .D(n65627), .S0(n65860), 
        .S1(n65756), .Q(n62223) );
  IMUX40 U68871 ( .A(n65620), .B(n65621), .C(n65622), .D(n65623), .S0(n65861), 
        .S1(n65756), .Q(n62221) );
  IMUX40 U68710 ( .A(n62220), .B(n62221), .C(n62222), .D(n62223), .S0(N1240), 
        .S1(n65918), .Q(n62219) );
  IMUX40 U9077 ( .A(n65724), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(n65727), 
        .S0(n65810), .S1(N704), .Q(n5275) );
  IMUX40 U9074 ( .A(n65736), .B(\GFill[13][0] ), .C(\GFill[14][0] ), .D(n65739), .S0(n65811), .S1(N704), .Q(n5278) );
  IMUX40 U9075 ( .A(n65732), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(n65735), 
        .S0(n65810), .S1(N704), .Q(n5276) );
  IMUX40 U8905 ( .A(n5275), .B(n5276), .C(n5277), .D(n5278), .S0(N706), .S1(
        N705), .Q(n5274) );
  IMUX40 U9073 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(n65710), .D(
        \GFill[19][0] ), .S0(n65811), .S1(N704), .Q(n5270) );
  IMUX40 U9070 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(n65722), .D(
        \GFill[31][0] ), .S0(n65811), .S1(N704), .Q(n5273) );
  IMUX40 U9071 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(n65718), .D(
        \GFill[27][0] ), .S0(n65811), .S1(N704), .Q(n5271) );
  IMUX40 U8904 ( .A(n5270), .B(n5271), .C(n5272), .D(n5273), .S0(N706), .S1(
        N705), .Q(n5269) );
  IMUX40 U10421 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65817), .S1(N716), .Q(n6555) );
  IMUX40 U10418 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65818), .S1(N716), .Q(n6558) );
  IMUX40 U10419 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65818), .S1(N716), .Q(n6556) );
  IMUX40 U10249 ( .A(n6555), .B(n6556), .C(n6557), .D(n6558), .S0(N718), .S1(
        N717), .Q(n6554) );
  IMUX40 U10417 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65818), .S1(N716), .Q(n6550) );
  IMUX40 U10414 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65818), .S1(N716), .Q(n6553) );
  IMUX40 U10415 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65818), .S1(N716), .Q(n6551) );
  IMUX40 U10248 ( .A(n6550), .B(n6551), .C(n6552), .D(n6553), .S0(N718), .S1(
        N717), .Q(n6549) );
  IMUX40 U11093 ( .A(n65724), .B(n65725), .C(\GFill[2][0] ), .D(n65727), .S0(
        n65820), .S1(N722), .Q(n7195) );
  IMUX40 U11090 ( .A(n65736), .B(n65737), .C(\GFill[14][0] ), .D(n65739), .S0(
        n65831), .S1(N722), .Q(n7198) );
  IMUX40 U11091 ( .A(n65732), .B(n65733), .C(\GFill[10][0] ), .D(n65735), .S0(
        n65831), .S1(N722), .Q(n7196) );
  IMUX40 U10921 ( .A(n7195), .B(n7196), .C(n7197), .D(n7198), .S0(N724), .S1(
        N723), .Q(n7194) );
  IMUX40 U11089 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(n65710), .D(
        \GFill[19][0] ), .S0(n65831), .S1(N722), .Q(n7190) );
  IMUX40 U11086 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(n65722), .D(
        \GFill[31][0] ), .S0(n65831), .S1(N722), .Q(n7193) );
  IMUX40 U11087 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(n65718), .D(
        \GFill[27][0] ), .S0(n65831), .S1(N722), .Q(n7191) );
  IMUX40 U10920 ( .A(n7190), .B(n7191), .C(n7192), .D(n7193), .S0(N724), .S1(
        N723), .Q(n7189) );
  IMUX40 U13109 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65825), .S1(N740), .Q(n9115) );
  IMUX40 U13106 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65824), .S1(N740), .Q(n9118) );
  IMUX40 U13107 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65824), .S1(N740), .Q(n9116) );
  IMUX40 U12937 ( .A(n9115), .B(n9116), .C(n9117), .D(n9118), .S0(N742), .S1(
        N741), .Q(n9114) );
  IMUX40 U13105 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65824), .S1(N740), .Q(n9110) );
  IMUX40 U13102 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65824), .S1(N740), .Q(n9113) );
  IMUX40 U13103 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65824), .S1(N740), .Q(n9111) );
  IMUX40 U12936 ( .A(n9110), .B(n9111), .C(n9112), .D(n9113), .S0(N742), .S1(
        N741), .Q(n9109) );
  IMUX40 U40661 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65813), .S1(N980), .Q(n35355) );
  IMUX40 U40658 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(n65674), .D(
        \OFill[15][0] ), .S0(n65813), .S1(N980), .Q(n35358) );
  IMUX40 U40659 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65813), .S1(N980), .Q(n35356) );
  IMUX40 U40489 ( .A(n35355), .B(n35356), .C(n35357), .D(n35358), .S0(N988), 
        .S1(N987), .Q(n35354) );
  IMUX40 U40657 ( .A(\OFill[16][0] ), .B(n65645), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65813), .S1(N980), .Q(n35350) );
  IMUX40 U40654 ( .A(\OFill[28][0] ), .B(n65657), .C(n65658), .D(
        \OFill[31][0] ), .S0(n65814), .S1(N980), .Q(n35353) );
  IMUX40 U40655 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(n65654), .D(
        n65655), .S0(n65814), .S1(N980), .Q(n35351) );
  IMUX40 U40488 ( .A(n35350), .B(n35351), .C(n35352), .D(n35353), .S0(N988), 
        .S1(N987), .Q(n35349) );
  IMUX40 U39989 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65791), .S1(n65924), .Q(n34715) );
  IMUX40 U39986 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65798), .S1(N1010), .Q(n34718) );
  IMUX40 U39987 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65802), .S1(N980), .Q(n34716) );
  IMUX40 U39817 ( .A(n34715), .B(n34716), .C(n34717), .D(n34718), .S0(N982), 
        .S1(N981), .Q(n34714) );
  IMUX40 U39985 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65806), .S1(n65924), .Q(n34710) );
  IMUX40 U39982 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65801), .S1(N980), .Q(n34713) );
  IMUX40 U39983 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65799), .S1(n65925), .Q(n34711) );
  IMUX40 U39816 ( .A(n34710), .B(n34711), .C(n34712), .D(n34713), .S0(N982), 
        .S1(N981), .Q(n34709) );
  IMUX40 U41333 ( .A(n65660), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(n65663), 
        .S0(n65815), .S1(N1004), .Q(n35995) );
  IMUX40 U41330 ( .A(n65672), .B(\OFill[13][0] ), .C(n65674), .D(n65675), .S0(
        n65815), .S1(N1004), .Q(n35998) );
  IMUX40 U41331 ( .A(n65668), .B(\OFill[9][0] ), .C(\OFill[10][0] ), .D(n65671), .S0(n65815), .S1(N1004), .Q(n35996) );
  IMUX40 U41161 ( .A(n35995), .B(n35996), .C(n35997), .D(n35998), .S0(N994), 
        .S1(N993), .Q(n35994) );
  IMUX40 U41329 ( .A(\OFill[16][0] ), .B(n65645), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65816), .S1(N1004), .Q(n35990) );
  IMUX40 U41326 ( .A(\OFill[28][0] ), .B(n65657), .C(n65658), .D(
        \OFill[31][0] ), .S0(n65816), .S1(N1004), .Q(n35993) );
  IMUX40 U41327 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(n65654), .D(
        n65655), .S0(n65816), .S1(N1004), .Q(n35991) );
  IMUX40 U41160 ( .A(n35990), .B(n35991), .C(n35992), .D(n35993), .S0(N994), 
        .S1(N993), .Q(n35989) );
  IMUX40 U42677 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65830), .S1(N716), .Q(n37275) );
  IMUX40 U42674 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65829), .S1(n65928), .Q(n37278) );
  IMUX40 U42675 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65829), .S1(N1004), .Q(n37276) );
  IMUX40 U42505 ( .A(n37275), .B(n37276), .C(n37277), .D(n37278), .S0(N1006), 
        .S1(N1005), .Q(n37274) );
  IMUX40 U42673 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65829), .S1(n65928), .Q(n37270) );
  IMUX40 U42670 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65828), .S1(N1004), .Q(n37273) );
  IMUX40 U42671 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65829), .S1(n65929), .Q(n37271) );
  IMUX40 U42504 ( .A(n37270), .B(n37271), .C(n37272), .D(n37273), .S0(N1006), 
        .S1(N1005), .Q(n37269) );
  IMUX40 U43349 ( .A(n65660), .B(\OFill[1][0] ), .C(n65662), .D(n65663), .S0(
        n65827), .S1(N1010), .Q(n37915) );
  IMUX40 U43346 ( .A(n65672), .B(\OFill[13][0] ), .C(\OFill[14][0] ), .D(
        n65675), .S0(n65827), .S1(n65924), .Q(n37918) );
  IMUX40 U43347 ( .A(n65668), .B(\OFill[9][0] ), .C(n65670), .D(n65671), .S0(
        n65827), .S1(n65925), .Q(n37916) );
  IMUX40 U43177 ( .A(n37915), .B(n37916), .C(n37917), .D(n37918), .S0(N1012), 
        .S1(N1011), .Q(n37914) );
  IMUX40 U43345 ( .A(\OFill[16][0] ), .B(n65645), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65827), .S1(N1010), .Q(n37910) );
  IMUX40 U43342 ( .A(\OFill[28][0] ), .B(n65657), .C(\OFill[30][0] ), .D(
        \OFill[31][0] ), .S0(n65826), .S1(n65925), .Q(n37913) );
  IMUX40 U43343 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(n65654), .D(
        n65655), .S0(n65826), .S1(N980), .Q(n37911) );
  IMUX40 U43176 ( .A(n37910), .B(n37911), .C(n37912), .D(n37913), .S0(N1012), 
        .S1(N1011), .Q(n37909) );
  IMUX40 U45365 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65822), .S1(N704), .Q(n39835) );
  IMUX40 U45362 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65822), .S1(n65926), .Q(n39838) );
  IMUX40 U45363 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65822), .S1(N1040), .Q(n39836) );
  IMUX40 U45193 ( .A(n39835), .B(n39836), .C(n39837), .D(n39838), .S0(N1030), 
        .S1(N1029), .Q(n39834) );
  IMUX40 U45361 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65822), .S1(n65927), .Q(n39830) );
  IMUX40 U45358 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(n65658), .D(
        \OFill[31][0] ), .S0(n65821), .S1(n65926), .Q(n39833) );
  IMUX40 U45359 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65822), .S1(n65927), .Q(n39831) );
  IMUX40 U45192 ( .A(n39830), .B(n39831), .C(n39832), .D(n39833), .S0(N1030), 
        .S1(N1029), .Q(n39829) );
  IMUX40 U27893 ( .A(n65724), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(n65727), 
        .S0(n65882), .S1(n65778), .Q(n23195) );
  IMUX40 U27890 ( .A(n65736), .B(\GFill[13][0] ), .C(\GFill[14][0] ), .D(
        n65739), .S0(n65880), .S1(n65774), .Q(n23198) );
  IMUX40 U27891 ( .A(n65732), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(n65735), .S0(n65881), .S1(n65778), .Q(n23196) );
  IMUX40 U27721 ( .A(n23195), .B(n23196), .C(n23197), .D(n23198), .S0(N874), 
        .S1(N873), .Q(n23194) );
  IMUX40 U27889 ( .A(n65708), .B(n65709), .C(\GFill[18][0] ), .D(n65711), .S0(
        n65876), .S1(n65762), .Q(n23190) );
  IMUX40 U27886 ( .A(n65720), .B(n65721), .C(\GFill[30][0] ), .D(n65723), .S0(
        n65869), .S1(n65772), .Q(n23193) );
  IMUX40 U27887 ( .A(n65716), .B(n65717), .C(\GFill[26][0] ), .D(n65719), .S0(
        n65907), .S1(n65760), .Q(n23191) );
  IMUX40 U27720 ( .A(n23190), .B(n23191), .C(n23192), .D(n23193), .S0(N874), 
        .S1(N873), .Q(n23189) );
  IMUX40 U26549 ( .A(n65724), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65793), .S1(n65534), .Q(n21915) );
  IMUX40 U26546 ( .A(n65736), .B(\GFill[13][0] ), .C(\GFill[14][0] ), .D(
        \GFill[15][0] ), .S0(n65792), .S1(n65534), .Q(n21918) );
  IMUX40 U26547 ( .A(n65732), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(
        \GFill[11][0] ), .S0(n65794), .S1(n65534), .Q(n21916) );
  IMUX40 U26377 ( .A(n21915), .B(n21916), .C(n21917), .D(n21918), .S0(N862), 
        .S1(N861), .Q(n21914) );
  IMUX40 U26545 ( .A(n65708), .B(\GFill[17][0] ), .C(\GFill[18][0] ), .D(
        \GFill[19][0] ), .S0(n65784), .S1(n65534), .Q(n21910) );
  IMUX40 U26542 ( .A(n65720), .B(\GFill[29][0] ), .C(\GFill[30][0] ), .D(
        \GFill[31][0] ), .S0(n65787), .S1(n65534), .Q(n21913) );
  IMUX40 U26543 ( .A(n65716), .B(\GFill[25][0] ), .C(\GFill[26][0] ), .D(
        \GFill[27][0] ), .S0(n65790), .S1(n65534), .Q(n21911) );
  IMUX40 U26376 ( .A(n21910), .B(n21911), .C(n21912), .D(n21913), .S0(N862), 
        .S1(N861), .Q(n21909) );
  IMUX40 U25877 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(n65726), .D(
        \GFill[3][0] ), .S0(N1207), .S1(n65773), .Q(n21275) );
  IMUX40 U25874 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(n65738), .D(
        \GFill[15][0] ), .S0(n65892), .S1(n65776), .Q(n21278) );
  IMUX40 U25875 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(n65734), .D(
        \GFill[11][0] ), .S0(n65869), .S1(n65778), .Q(n21276) );
  IMUX40 U25705 ( .A(n21275), .B(n21276), .C(n21277), .D(n21278), .S0(N856), 
        .S1(N855), .Q(n21274) );
  IMUX40 U25873 ( .A(\GFill[16][0] ), .B(n65709), .C(\GFill[18][0] ), .D(
        \GFill[19][0] ), .S0(n65873), .S1(n65777), .Q(n21270) );
  IMUX40 U25870 ( .A(\GFill[28][0] ), .B(n65721), .C(\GFill[30][0] ), .D(
        \GFill[31][0] ), .S0(n65884), .S1(n65776), .Q(n21273) );
  IMUX40 U25871 ( .A(\GFill[24][0] ), .B(n65717), .C(\GFill[26][0] ), .D(
        \GFill[27][0] ), .S0(n65899), .S1(n65763), .Q(n21271) );
  IMUX40 U25704 ( .A(n21270), .B(n21271), .C(n21272), .D(n21273), .S0(N856), 
        .S1(N855), .Q(n21269) );
  IMUX40 U60149 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65886), .S1(n65765), .Q(n53915) );
  IMUX40 U60146 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65878), .S1(n65771), .Q(n53918) );
  IMUX40 U60147 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65859), .S1(n65763), .Q(n53916) );
  IMUX40 U59977 ( .A(n53915), .B(n53916), .C(n53917), .D(n53918), .S0(N1162), 
        .S1(N1161), .Q(n53914) );
  IMUX40 U60145 ( .A(n65644), .B(\OFill[17][0] ), .C(n65646), .D(n65647), .S0(
        n65849), .S1(n65771), .Q(n53910) );
  IMUX40 U60142 ( .A(n65656), .B(\OFill[29][0] ), .C(\OFill[30][0] ), .D(
        n65659), .S0(n65869), .S1(n65771), .Q(n53913) );
  IMUX40 U60143 ( .A(n65652), .B(n65653), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65862), .S1(n65771), .Q(n53911) );
  IMUX40 U59976 ( .A(n53910), .B(n53911), .C(n53912), .D(n53913), .S0(N1162), 
        .S1(N1161), .Q(n53909) );
  IMUX40 U58805 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(n65662), .D(n65663), 
        .S0(n65818), .S1(n65537), .Q(n52635) );
  IMUX40 U58802 ( .A(n65672), .B(n65673), .C(\OFill[14][0] ), .D(n65675), .S0(
        n65825), .S1(n65537), .Q(n52638) );
  IMUX40 U58803 ( .A(n65668), .B(\OFill[9][0] ), .C(n65670), .D(n65671), .S0(
        n65826), .S1(n65537), .Q(n52636) );
  IMUX40 U58633 ( .A(n52635), .B(n52636), .C(n52637), .D(n52638), .S0(N1150), 
        .S1(N1149), .Q(n52634) );
  IMUX40 U58801 ( .A(n65644), .B(\OFill[17][0] ), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65822), .S1(n65537), .Q(n52630) );
  IMUX40 U58798 ( .A(n65656), .B(\OFill[29][0] ), .C(\OFill[30][0] ), .D(
        \OFill[31][0] ), .S0(n65823), .S1(n65537), .Q(n52633) );
  IMUX40 U58799 ( .A(n65652), .B(\OFill[25][0] ), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65824), .S1(n65537), .Q(n52631) );
  IMUX40 U58632 ( .A(n52630), .B(n52631), .C(n52632), .D(n52633), .S0(N1150), 
        .S1(N1149), .Q(n52629) );
  IMUX40 U58133 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65887), .S1(n65759), .Q(n51995) );
  IMUX40 U58130 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65876), .S1(n65773), .Q(n51998) );
  IMUX40 U58131 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65905), .S1(n65781), .Q(n51996) );
  IMUX40 U57961 ( .A(n51995), .B(n51996), .C(n51997), .D(n51998), .S0(N1144), 
        .S1(N1143), .Q(n51994) );
  IMUX40 U58129 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65836), .S1(n65780), .Q(n51990) );
  IMUX40 U58126 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65852), .S1(n65773), .Q(n51993) );
  IMUX40 U58127 ( .A(\OFill[24][0] ), .B(n65653), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65878), .S1(n65781), .Q(n51991) );
  IMUX40 U57960 ( .A(n51990), .B(n51991), .C(n51992), .D(n51993), .S0(N1144), 
        .S1(N1143), .Q(n51989) );
  IMUX40 U56789 ( .A(n65660), .B(n65661), .C(\OFill[2][0] ), .D(\OFill[3][0] ), 
        .S0(n65783), .S1(n65538), .Q(n50715) );
  IMUX40 U56786 ( .A(n65672), .B(\OFill[13][0] ), .C(\OFill[14][0] ), .D(
        \OFill[15][0] ), .S0(n65784), .S1(n65538), .Q(n50718) );
  IMUX40 U56787 ( .A(n65668), .B(n65669), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65783), .S1(n65538), .Q(n50716) );
  IMUX40 U56617 ( .A(n50715), .B(n50716), .C(n50717), .D(n50718), .S0(N1132), 
        .S1(N1131), .Q(n50714) );
  IMUX40 U56785 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65784), 
        .S1(n65538), .Q(n50710) );
  IMUX40 U56782 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65784), 
        .S1(n65538), .Q(n50713) );
  IMUX40 U56783 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65784), 
        .S1(n65538), .Q(n50711) );
  IMUX40 U56616 ( .A(n50710), .B(n50711), .C(n50712), .D(n50713), .S0(N1132), 
        .S1(N1131), .Q(n50709) );
  IMUX40 U56117 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65862), .S1(n65778), .Q(n50075) );
  IMUX40 U56114 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65880), .S1(n65769), .Q(n50078) );
  IMUX40 U56115 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65882), .S1(n65762), .Q(n50076) );
  IMUX40 U55945 ( .A(n50075), .B(n50076), .C(n50077), .D(n50078), .S0(N1126), 
        .S1(N1125), .Q(n50074) );
  IMUX40 U56113 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65879), .S1(n65777), .Q(n50070) );
  IMUX40 U56110 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65879), .S1(n65759), .Q(n50073) );
  IMUX40 U56111 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65898), .S1(n65780), .Q(n50071) );
  IMUX40 U55944 ( .A(n50070), .B(n50071), .C(n50072), .D(n50073), .S0(N1126), 
        .S1(N1125), .Q(n50069) );
  IMUX40 U57461 ( .A(n65660), .B(n65661), .C(\OFill[2][0] ), .D(\OFill[3][0] ), 
        .S0(n65883), .S1(n65748), .Q(n51355) );
  IMUX40 U57458 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65835), .S1(n65748), .Q(n51358) );
  IMUX40 U57459 ( .A(\OFill[8][0] ), .B(n65669), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65899), .S1(n65748), .Q(n51356) );
  IMUX40 U57289 ( .A(n51355), .B(n51356), .C(n51357), .D(n51358), .S0(N1138), 
        .S1(n65919), .Q(n51354) );
  IMUX40 U57457 ( .A(n65644), .B(\OFill[17][0] ), .C(n65646), .D(n65647), .S0(
        n65835), .S1(n65748), .Q(n51350) );
  IMUX40 U57454 ( .A(n65656), .B(\OFill[29][0] ), .C(n65658), .D(n65659), .S0(
        n65857), .S1(n65748), .Q(n51353) );
  IMUX40 U57455 ( .A(n65652), .B(\OFill[25][0] ), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65836), .S1(n65748), .Q(n51351) );
  IMUX40 U57288 ( .A(n51350), .B(n51351), .C(n51352), .D(n51353), .S0(N1138), 
        .S1(n65919), .Q(n51349) );
  IMUX40 U39317 ( .A(n65724), .B(n65725), .C(n65726), .D(n65727), .S0(n65894), 
        .S1(n65769), .Q(n34075) );
  IMUX40 U39314 ( .A(n65736), .B(n65737), .C(n65738), .D(n65739), .S0(n65906), 
        .S1(n65769), .Q(n34078) );
  IMUX40 U39315 ( .A(n65732), .B(n65733), .C(n65734), .D(n65735), .S0(n65890), 
        .S1(n65769), .Q(n34076) );
  IMUX40 U39145 ( .A(n34075), .B(n34076), .C(n34077), .D(n34078), .S0(N976), 
        .S1(N975), .Q(n34074) );
  IMUX40 U39313 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65900), 
        .S1(n65769), .Q(n34070) );
  IMUX40 U39310 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65865), 
        .S1(n65768), .Q(n34073) );
  IMUX40 U39311 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65891), 
        .S1(n65768), .Q(n34071) );
  IMUX40 U39144 ( .A(n34070), .B(n34071), .C(n34072), .D(n34073), .S0(N976), 
        .S1(N975), .Q(n34069) );
  IMUX40 U71573 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65906), 
        .S1(n65767), .Q(n64795) );
  IMUX40 U71570 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65850), 
        .S1(n65766), .Q(n64798) );
  IMUX40 U71571 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65862), 
        .S1(n65766), .Q(n64796) );
  IMUX40 U71401 ( .A(n64795), .B(n64796), .C(n64797), .D(n64798), .S0(N1264), 
        .S1(N1263), .Q(n64794) );
  IMUX40 U71569 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65859), 
        .S1(n65764), .Q(n64790) );
  IMUX40 U71566 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65834), 
        .S1(n65766), .Q(n64793) );
  IMUX40 U71567 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65897), 
        .S1(n65766), .Q(n64791) );
  IMUX40 U71400 ( .A(n64790), .B(n64791), .C(n64792), .D(n64793), .S0(N1264), 
        .S1(N1263), .Q(n64789) );
  IMUX40 U35285 ( .A(\GFill[0][0] ), .B(n65725), .C(n65726), .D(n65727), .S0(
        n65832), .S1(n65755), .Q(n30235) );
  IMUX40 U35282 ( .A(\GFill[12][0] ), .B(n65737), .C(n65738), .D(n65739), .S0(
        n65856), .S1(n65755), .Q(n30238) );
  IMUX40 U35283 ( .A(\GFill[8][0] ), .B(n65733), .C(n65734), .D(n65735), .S0(
        n65895), .S1(n65755), .Q(n30236) );
  IMUX40 U35113 ( .A(n30235), .B(n30236), .C(n30237), .D(n30238), .S0(N940), 
        .S1(n65918), .Q(n30234) );
  IMUX40 U35281 ( .A(\GFill[16][0] ), .B(n65709), .C(n65710), .D(n65711), .S0(
        n65874), .S1(n65755), .Q(n30230) );
  IMUX40 U35278 ( .A(\GFill[28][0] ), .B(n65721), .C(n65722), .D(n65723), .S0(
        n65841), .S1(n65754), .Q(n30233) );
  IMUX40 U35279 ( .A(\GFill[24][0] ), .B(n65717), .C(n65718), .D(n65719), .S0(
        n65868), .S1(n65754), .Q(n30231) );
  IMUX40 U35112 ( .A(n30230), .B(n30231), .C(n30232), .D(n30233), .S0(N940), 
        .S1(n65918), .Q(n30229) );
  IMUX40 U67541 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65840), 
        .S1(n65746), .Q(n60955) );
  IMUX40 U67538 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65870), 
        .S1(n65747), .Q(n60958) );
  IMUX40 U67539 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65895), 
        .S1(n65747), .Q(n60956) );
  IMUX40 U67369 ( .A(n60955), .B(n60956), .C(n60957), .D(n60958), .S0(N1228), 
        .S1(n65917), .Q(n60954) );
  IMUX40 U67537 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65868), 
        .S1(n65747), .Q(n60950) );
  IMUX40 U67534 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65908), 
        .S1(n65747), .Q(n60953) );
  IMUX40 U67535 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65887), 
        .S1(n65747), .Q(n60951) );
  IMUX40 U67368 ( .A(n60950), .B(n60951), .C(n60952), .D(n60953), .S0(N1228), 
        .S1(n65917), .Q(n60949) );
  IMUX40 U37973 ( .A(n65724), .B(n65725), .C(n65726), .D(n65727), .S0(n65868), 
        .S1(n65753), .Q(n32795) );
  IMUX40 U37970 ( .A(n65736), .B(n65737), .C(n65738), .D(n65739), .S0(n65847), 
        .S1(n65751), .Q(n32798) );
  IMUX40 U37971 ( .A(n65732), .B(n65733), .C(n65734), .D(n65735), .S0(n65858), 
        .S1(n65753), .Q(n32796) );
  IMUX40 U37801 ( .A(n32795), .B(n32796), .C(n32797), .D(n32798), .S0(N964), 
        .S1(n65916), .Q(n32794) );
  IMUX40 U37969 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65882), 
        .S1(n65748), .Q(n32790) );
  IMUX40 U37966 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65888), 
        .S1(n65747), .Q(n32793) );
  IMUX40 U37967 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65861), 
        .S1(n65750), .Q(n32791) );
  IMUX40 U37800 ( .A(n32790), .B(n32791), .C(n32792), .D(n32793), .S0(N964), 
        .S1(n65918), .Q(n32789) );
  IMUX40 U36629 ( .A(n65724), .B(n65725), .C(n65726), .D(n65727), .S0(n65870), 
        .S1(n65756), .Q(n31515) );
  IMUX40 U36626 ( .A(n65736), .B(n65737), .C(n65738), .D(n65739), .S0(n65855), 
        .S1(n65756), .Q(n31518) );
  IMUX40 U36627 ( .A(n65732), .B(n65733), .C(n65734), .D(n65735), .S0(n65844), 
        .S1(n65756), .Q(n31516) );
  IMUX40 U36457 ( .A(n31515), .B(n31516), .C(n31517), .D(n31518), .S0(N952), 
        .S1(n65918), .Q(n31514) );
  IMUX40 U36625 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65907), 
        .S1(n65756), .Q(n31510) );
  IMUX40 U36622 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65875), 
        .S1(n65755), .Q(n31513) );
  IMUX40 U36623 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65881), 
        .S1(n65755), .Q(n31511) );
  IMUX40 U36456 ( .A(n31510), .B(n31511), .C(n31512), .D(n31513), .S0(N952), 
        .S1(n65916), .Q(n31509) );
  IMUX40 U70229 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65832), 
        .S1(n65754), .Q(n63515) );
  IMUX40 U70226 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65864), 
        .S1(n65752), .Q(n63518) );
  IMUX40 U70227 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65841), 
        .S1(n65749), .Q(n63516) );
  IMUX40 U70057 ( .A(n63515), .B(n63516), .C(n63517), .D(n63518), .S0(N1252), 
        .S1(n65916), .Q(n63514) );
  IMUX40 U70225 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65898), 
        .S1(n65746), .Q(n63510) );
  IMUX40 U70222 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65859), 
        .S1(N1208), .Q(n63513) );
  IMUX40 U70223 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65840), 
        .S1(n65755), .Q(n63511) );
  IMUX40 U70056 ( .A(n63510), .B(n63511), .C(n63512), .D(n63513), .S0(N1252), 
        .S1(n65916), .Q(n63509) );
  IMUX40 U68885 ( .A(n65660), .B(n65661), .C(n65662), .D(n65663), .S0(n65879), 
        .S1(n65757), .Q(n62235) );
  IMUX40 U68882 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65885), 
        .S1(n65757), .Q(n62238) );
  IMUX40 U68883 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65835), 
        .S1(n65757), .Q(n62236) );
  IMUX40 U68713 ( .A(n62235), .B(n62236), .C(n62237), .D(n62238), .S0(N1240), 
        .S1(n65918), .Q(n62234) );
  IMUX40 U68881 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65909), 
        .S1(n65757), .Q(n62230) );
  IMUX40 U68878 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65842), 
        .S1(n65757), .Q(n62233) );
  IMUX40 U68879 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65905), 
        .S1(n65757), .Q(n62231) );
  IMUX40 U68712 ( .A(n62230), .B(n62231), .C(n62232), .D(n62233), .S0(N1240), 
        .S1(n65916), .Q(n62229) );
  IMUX40 U48717 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65818), .S1(n65912), .Q(n43025) );
  IMUX40 U48714 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65809), .S1(N1082), .Q(n43028) );
  IMUX40 U48715 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65808), .S1(n65922), .Q(n43026) );
  IMUX40 U48551 ( .A(n43025), .B(n43026), .C(n43027), .D(n43028), .S0(N1060), 
        .S1(N1059), .Q(n43024) );
  IMUX40 U48713 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65783), .S1(n65911), .Q(n43020) );
  IMUX40 U48710 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65827), .S1(n65537), .Q(n43023) );
  IMUX40 U48711 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65800), .S1(n65537), .Q(n43021) );
  IMUX40 U48550 ( .A(n43020), .B(n43021), .C(n43022), .D(n43023), .S0(N1060), 
        .S1(N1059), .Q(n43019) );
  IMUX40 U48045 ( .A(n65628), .B(\OFill[33][0] ), .C(\OFill[34][0] ), .D(
        \OFill[35][0] ), .S0(n65866), .S1(n65781), .Q(n42385) );
  IMUX40 U48042 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65865), .S1(n65775), .Q(n42388) );
  IMUX40 U48043 ( .A(n65636), .B(\OFill[41][0] ), .C(\OFill[42][0] ), .D(
        \OFill[43][0] ), .S0(n65866), .S1(n65776), .Q(n42386) );
  IMUX40 U47879 ( .A(n42385), .B(n42386), .C(n42387), .D(n42388), .S0(N1054), 
        .S1(N1053), .Q(n42384) );
  IMUX40 U48041 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65865), .S1(n65774), .Q(n42380) );
  IMUX40 U48038 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65864), .S1(n65767), .Q(n42383) );
  IMUX40 U48039 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65864), .S1(n65773), .Q(n42381) );
  IMUX40 U47878 ( .A(n42380), .B(n42381), .C(n42382), .D(n42383), .S0(N1054), 
        .S1(N1053), .Q(n42379) );
  IMUX40 U50733 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65873), .S1(n65776), .Q(n44945) );
  IMUX40 U50730 ( .A(n65640), .B(\OFill[45][0] ), .C(\OFill[46][0] ), .D(
        \OFill[47][0] ), .S0(n65834), .S1(n65781), .Q(n44948) );
  IMUX40 U50731 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65874), .S1(n65777), .Q(n44946) );
  IMUX40 U50567 ( .A(n44945), .B(n44946), .C(n44947), .D(n44948), .S0(N1078), 
        .S1(N1077), .Q(n44944) );
  IMUX40 U50729 ( .A(n65612), .B(\OFill[49][0] ), .C(\OFill[50][0] ), .D(
        \OFill[51][0] ), .S0(n65897), .S1(n65775), .Q(n44940) );
  IMUX40 U50726 ( .A(n65624), .B(\OFill[61][0] ), .C(\OFill[62][0] ), .D(
        \OFill[63][0] ), .S0(n65874), .S1(n65767), .Q(n44943) );
  IMUX40 U50727 ( .A(n65620), .B(\OFill[57][0] ), .C(\OFill[58][0] ), .D(
        \OFill[59][0] ), .S0(n65872), .S1(n65764), .Q(n44941) );
  IMUX40 U50566 ( .A(n44940), .B(n44941), .C(n44942), .D(n44943), .S0(N1078), 
        .S1(N1077), .Q(n44939) );
  IMUX40 U64845 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(n65630), .D(
        \OFill[35][0] ), .S0(n65803), .S1(n65912), .Q(n58385) );
  IMUX40 U64842 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(n65642), .D(
        \OFill[47][0] ), .S0(n65799), .S1(N1082), .Q(n58388) );
  IMUX40 U64843 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(n65638), .D(
        \OFill[43][0] ), .S0(n65800), .S1(n65537), .Q(n58386) );
  IMUX40 U64679 ( .A(n58385), .B(n58386), .C(n58387), .D(n58388), .S0(N1204), 
        .S1(N1203), .Q(n58384) );
  IMUX40 U64841 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(n65614), .D(
        \OFill[51][0] ), .S0(n65830), .S1(n65912), .Q(n58380) );
  IMUX40 U64838 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(n65626), .D(
        \OFill[63][0] ), .S0(n65820), .S1(n65923), .Q(n58383) );
  IMUX40 U64839 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(n65622), .D(
        \OFill[59][0] ), .S0(n65785), .S1(n65923), .Q(n58381) );
  IMUX40 U64678 ( .A(n58380), .B(n58381), .C(n58382), .D(n58383), .S0(N1204), 
        .S1(N1203), .Q(n58379) );
  IMUX40 U15789 ( .A(n65692), .B(\GFill[33][0] ), .C(\GFill[34][0] ), .D(
        \GFill[35][0] ), .S0(n65861), .S1(n65763), .Q(n11665) );
  IMUX40 U15786 ( .A(n65704), .B(\GFill[45][0] ), .C(\GFill[46][0] ), .D(
        \GFill[47][0] ), .S0(n65862), .S1(n65769), .Q(n11668) );
  IMUX40 U15787 ( .A(n65700), .B(\GFill[41][0] ), .C(\GFill[42][0] ), .D(
        \GFill[43][0] ), .S0(n65862), .S1(n65760), .Q(n11666) );
  IMUX40 U15623 ( .A(n11665), .B(n11666), .C(n11667), .D(n11668), .S0(N1054), 
        .S1(N1053), .Q(n11664) );
  IMUX40 U15785 ( .A(n65676), .B(\GFill[49][0] ), .C(\GFill[50][0] ), .D(
        \GFill[51][0] ), .S0(n65863), .S1(n65781), .Q(n11660) );
  IMUX40 U15782 ( .A(n65688), .B(\GFill[61][0] ), .C(\GFill[62][0] ), .D(
        \GFill[63][0] ), .S0(n65864), .S1(n65759), .Q(n11663) );
  IMUX40 U15783 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65863), .S1(n65780), .Q(n11661) );
  IMUX40 U15622 ( .A(n11660), .B(n11661), .C(n11662), .D(n11663), .S0(N1054), 
        .S1(N1053), .Q(n11659) );
  IMUX40 U34605 ( .A(\GFill[32][0] ), .B(n65693), .C(n65694), .D(n65695), .S0(
        n65808), .S1(N860), .Q(n29585) );
  IMUX40 U34602 ( .A(\GFill[44][0] ), .B(n65705), .C(n65706), .D(n65707), .S0(
        n65821), .S1(N1082), .Q(n29588) );
  IMUX40 U34603 ( .A(\GFill[40][0] ), .B(n65701), .C(n65702), .D(n65703), .S0(
        n65803), .S1(n65923), .Q(n29586) );
  IMUX40 U34439 ( .A(n29585), .B(n29586), .C(n29587), .D(n29588), .S0(N1222), 
        .S1(N1221), .Q(n29584) );
  IMUX40 U34601 ( .A(\GFill[48][0] ), .B(n65677), .C(n65678), .D(n65679), .S0(
        n65799), .S1(N1082), .Q(n29580) );
  IMUX40 U34598 ( .A(\GFill[60][0] ), .B(n65689), .C(n65690), .D(n65691), .S0(
        n65798), .S1(N1130), .Q(n29583) );
  IMUX40 U34599 ( .A(\GFill[56][0] ), .B(n65685), .C(n65686), .D(n65687), .S0(
        n65802), .S1(N1148), .Q(n29581) );
  IMUX40 U34438 ( .A(n29580), .B(n29581), .C(n29582), .D(n29583), .S0(N1222), 
        .S1(N1221), .Q(n29579) );
  IMUX40 U33933 ( .A(\GFill[32][0] ), .B(n65693), .C(n65694), .D(n65695), .S0(
        n65877), .S1(n65760), .Q(n28945) );
  IMUX40 U33930 ( .A(\GFill[44][0] ), .B(n65705), .C(n65706), .D(n65707), .S0(
        n65840), .S1(n65761), .Q(n28948) );
  IMUX40 U33931 ( .A(\GFill[40][0] ), .B(n65701), .C(n65702), .D(n65703), .S0(
        n65871), .S1(n65761), .Q(n28946) );
  IMUX40 U33767 ( .A(n28945), .B(n28946), .C(n28947), .D(n28948), .S0(N1216), 
        .S1(N1215), .Q(n28944) );
  IMUX40 U33929 ( .A(\GFill[48][0] ), .B(n65677), .C(n65678), .D(n65679), .S0(
        n65897), .S1(n65761), .Q(n28940) );
  IMUX40 U33926 ( .A(\GFill[60][0] ), .B(n65689), .C(n65690), .D(n65691), .S0(
        n65904), .S1(n65762), .Q(n28943) );
  IMUX40 U33927 ( .A(\GFill[56][0] ), .B(n65685), .C(n65686), .D(n65687), .S0(
        n65886), .S1(n65761), .Q(n28941) );
  IMUX40 U33766 ( .A(n28940), .B(n28941), .C(n28942), .D(n28943), .S0(N1216), 
        .S1(N1215), .Q(n28939) );
  IMUX40 U66861 ( .A(\OFill[32][0] ), .B(n65629), .C(n65630), .D(n65631), .S0(
        n65814), .S1(N1220), .Q(n60305) );
  IMUX40 U66858 ( .A(\OFill[44][0] ), .B(n65641), .C(n65642), .D(n65643), .S0(
        n65826), .S1(n65923), .Q(n60308) );
  IMUX40 U66859 ( .A(\OFill[40][0] ), .B(n65637), .C(n65638), .D(n65639), .S0(
        n65830), .S1(N1130), .Q(n60306) );
  IMUX40 U66695 ( .A(n60305), .B(n60306), .C(n60307), .D(n60308), .S0(N1222), 
        .S1(N1221), .Q(n60304) );
  IMUX40 U66857 ( .A(\OFill[48][0] ), .B(n65613), .C(n65614), .D(n65615), .S0(
        n65823), .S1(n65743), .Q(n60300) );
  IMUX40 U66854 ( .A(\OFill[60][0] ), .B(n65625), .C(n65626), .D(n65627), .S0(
        n65824), .S1(n65911), .Q(n60303) );
  IMUX40 U66855 ( .A(\OFill[56][0] ), .B(n65621), .C(n65622), .D(n65623), .S0(
        n65825), .S1(n65743), .Q(n60301) );
  IMUX40 U66694 ( .A(n60300), .B(n60301), .C(n60302), .D(n60303), .S0(N1222), 
        .S1(N1221), .Q(n60299) );
  IMUX40 U66189 ( .A(\OFill[32][0] ), .B(n65629), .C(n65630), .D(n65631), .S0(
        n65838), .S1(n65763), .Q(n59665) );
  IMUX40 U66186 ( .A(\OFill[44][0] ), .B(n65641), .C(n65642), .D(n65643), .S0(
        n65838), .S1(n65762), .Q(n59668) );
  IMUX40 U66187 ( .A(\OFill[40][0] ), .B(n65637), .C(n65638), .D(n65639), .S0(
        n65857), .S1(n65763), .Q(n59666) );
  IMUX40 U66023 ( .A(n59665), .B(n59666), .C(n59667), .D(n59668), .S0(N1216), 
        .S1(N1215), .Q(n59664) );
  IMUX40 U66185 ( .A(\OFill[48][0] ), .B(n65613), .C(n65614), .D(n65615), .S0(
        n65884), .S1(n65762), .Q(n59660) );
  IMUX40 U66182 ( .A(\OFill[60][0] ), .B(n65625), .C(n65626), .D(n65627), .S0(
        n65865), .S1(n65762), .Q(n59663) );
  IMUX40 U66183 ( .A(\OFill[56][0] ), .B(n65621), .C(n65622), .D(n65623), .S0(
        n65907), .S1(n65762), .Q(n59661) );
  IMUX40 U66022 ( .A(n59660), .B(n59661), .C(n59662), .D(n59663), .S0(N1216), 
        .S1(N1215), .Q(n59659) );
  IMUX40 U21837 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65847), .S1(n65774), .Q(n17425) );
  IMUX40 U21834 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65848), .S1(n65766), .Q(n17428) );
  IMUX40 U21835 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65847), .S1(n65761), .Q(n17426) );
  IMUX40 U21671 ( .A(n17425), .B(n17426), .C(n17427), .D(n17428), .S0(N1108), 
        .S1(N1107), .Q(n17424) );
  IMUX40 U21833 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65848), .S1(n65773), .Q(n17420) );
  IMUX40 U21830 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65849), .S1(n65770), .Q(n17423) );
  IMUX40 U21831 ( .A(n65684), .B(\GFill[57][0] ), .C(\GFill[58][0] ), .D(
        \GFill[59][0] ), .S0(n65849), .S1(n65775), .Q(n17421) );
  IMUX40 U21670 ( .A(n17420), .B(n17421), .C(n17422), .D(n17423), .S0(N1108), 
        .S1(N1107), .Q(n17419) );
  IMUX40 U28557 ( .A(\GFill[32][0] ), .B(\GFill[33][0] ), .C(\GFill[34][0] ), 
        .D(\GFill[35][0] ), .S0(n65872), .S1(n65751), .Q(n23825) );
  IMUX40 U28554 ( .A(\GFill[44][0] ), .B(\GFill[45][0] ), .C(\GFill[46][0] ), 
        .D(\GFill[47][0] ), .S0(n65874), .S1(n65751), .Q(n23828) );
  IMUX40 U28555 ( .A(\GFill[40][0] ), .B(\GFill[41][0] ), .C(\GFill[42][0] ), 
        .D(\GFill[43][0] ), .S0(n65890), .S1(n65751), .Q(n23826) );
  IMUX40 U28391 ( .A(n23825), .B(n23826), .C(n23827), .D(n23828), .S0(N1168), 
        .S1(n65915), .Q(n23824) );
  IMUX40 U28553 ( .A(\GFill[48][0] ), .B(\GFill[49][0] ), .C(\GFill[50][0] ), 
        .D(\GFill[51][0] ), .S0(n65909), .S1(n65751), .Q(n23820) );
  IMUX40 U28550 ( .A(\GFill[60][0] ), .B(\GFill[61][0] ), .C(\GFill[62][0] ), 
        .D(\GFill[63][0] ), .S0(n65860), .S1(n65750), .Q(n23823) );
  IMUX40 U28551 ( .A(\GFill[56][0] ), .B(\GFill[57][0] ), .C(\GFill[58][0] ), 
        .D(\GFill[59][0] ), .S0(n65870), .S1(n65751), .Q(n23821) );
  IMUX40 U28390 ( .A(n23820), .B(n23821), .C(n23822), .D(n23823), .S0(N1168), 
        .S1(n65916), .Q(n23819) );
  IMUX40 U60813 ( .A(\OFill[32][0] ), .B(\OFill[33][0] ), .C(\OFill[34][0] ), 
        .D(\OFill[35][0] ), .S0(n65853), .S1(n65750), .Q(n54545) );
  IMUX40 U60810 ( .A(\OFill[44][0] ), .B(\OFill[45][0] ), .C(\OFill[46][0] ), 
        .D(\OFill[47][0] ), .S0(n65894), .S1(n65750), .Q(n54548) );
  IMUX40 U60811 ( .A(\OFill[40][0] ), .B(\OFill[41][0] ), .C(\OFill[42][0] ), 
        .D(\OFill[43][0] ), .S0(n65884), .S1(n65750), .Q(n54546) );
  IMUX40 U60647 ( .A(n54545), .B(n54546), .C(n54547), .D(n54548), .S0(N1168), 
        .S1(n65916), .Q(n54544) );
  IMUX40 U60809 ( .A(\OFill[48][0] ), .B(\OFill[49][0] ), .C(\OFill[50][0] ), 
        .D(\OFill[51][0] ), .S0(n65894), .S1(n65750), .Q(n54540) );
  IMUX40 U60806 ( .A(\OFill[60][0] ), .B(\OFill[61][0] ), .C(\OFill[62][0] ), 
        .D(\OFill[63][0] ), .S0(n65887), .S1(n65750), .Q(n54543) );
  IMUX40 U60807 ( .A(\OFill[56][0] ), .B(\OFill[57][0] ), .C(\OFill[58][0] ), 
        .D(\OFill[59][0] ), .S0(n65888), .S1(n65750), .Q(n54541) );
  IMUX40 U60646 ( .A(n54540), .B(n54541), .C(n54542), .D(n54543), .S0(N1168), 
        .S1(n65915), .Q(n54539) );
  IMUX40 U9745 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65798), .S1(N998), .Q(n5910) );
  IMUX40 U9742 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65811), .S1(n65935), .Q(n5913) );
  IMUX40 U9743 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65810), .S1(N998), .Q(n5911) );
  IMUX40 U9576 ( .A(n5910), .B(n5911), .C(n5912), .D(n5913), .S0(N1000), .S1(
        N999), .Q(n5909) );
  IMUX40 U12433 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65802), .S1(N1022), .Q(n8470) );
  IMUX40 U12430 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65802), .S1(n65933), .Q(n8473) );
  IMUX40 U12431 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65802), .S1(N1016), .Q(n8471) );
  IMUX40 U12264 ( .A(n8470), .B(n8471), .C(n8472), .D(n8473), .S0(N1024), .S1(
        N1023), .Q(n8469) );
  IMUX40 U11761 ( .A(n65708), .B(\GFill[17][0] ), .C(\GFill[18][0] ), .D(
        n65711), .S0(n65792), .S1(n65933), .Q(n7830) );
  IMUX40 U11758 ( .A(n65720), .B(\GFill[29][0] ), .C(\GFill[30][0] ), .D(
        n65723), .S0(n65782), .S1(n65933), .Q(n7833) );
  IMUX40 U11759 ( .A(n65716), .B(\GFill[25][0] ), .C(\GFill[26][0] ), .D(
        n65719), .S0(n65782), .S1(n65932), .Q(n7831) );
  IMUX40 U11592 ( .A(n7830), .B(n7831), .C(n7832), .D(n7833), .S0(N1018), .S1(
        N1017), .Q(n7829) );
  IMUX40 U13777 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65789), .S1(N1034), .Q(n9750) );
  IMUX40 U13774 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65792), .S1(n65929), .Q(n9753) );
  IMUX40 U13775 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65801), .S1(N1034), .Q(n9751) );
  IMUX40 U13608 ( .A(n9750), .B(n9751), .C(n9752), .D(n9753), .S0(N1036), .S1(
        N1035), .Q(n9749) );
  IMUX40 U15121 ( .A(n65708), .B(n65709), .C(\GFill[18][0] ), .D(n65711), .S0(
        n65794), .S1(N1046), .Q(n11030) );
  IMUX40 U15118 ( .A(n65720), .B(n65721), .C(\GFill[30][0] ), .D(n65723), .S0(
        n65794), .S1(N1010), .Q(n11033) );
  IMUX40 U15119 ( .A(n65716), .B(n65717), .C(\GFill[26][0] ), .D(n65719), .S0(
        n65794), .S1(n65925), .Q(n11031) );
  IMUX40 U14952 ( .A(n11030), .B(n11031), .C(n11032), .D(n11033), .S0(N1048), 
        .S1(N1047), .Q(n11029) );
  IMUX40 U14449 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65823), .S1(N1040), .Q(n10390) );
  IMUX40 U14446 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65824), .S1(n65927), .Q(n10393) );
  IMUX40 U14447 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65825), .S1(N1040), .Q(n10391) );
  IMUX40 U14280 ( .A(n10390), .B(n10391), .C(n10392), .D(n10393), .S0(N1042), 
        .S1(N1041), .Q(n10389) );
  IMUX40 U42001 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65801), .S1(n65934), .Q(n36630) );
  IMUX40 U41998 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(n65658), .D(
        \OFill[31][0] ), .S0(n65801), .S1(n65934), .Q(n36633) );
  IMUX40 U41999 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65801), .S1(n65934), .Q(n36631) );
  IMUX40 U41832 ( .A(n36630), .B(n36631), .C(n36632), .D(n36633), .S0(N1000), 
        .S1(N999), .Q(n36629) );
  IMUX40 U44689 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65805), .S1(n65932), .Q(n39190) );
  IMUX40 U44686 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65806), .S1(n65930), .Q(n39193) );
  IMUX40 U44687 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65806), .S1(n65933), .Q(n39191) );
  IMUX40 U44520 ( .A(n39190), .B(n39191), .C(n39192), .D(n39193), .S0(N1024), 
        .S1(N1023), .Q(n39189) );
  IMUX40 U44017 ( .A(n65644), .B(\OFill[17][0] ), .C(\OFill[18][0] ), .D(
        n65647), .S0(n65783), .S1(n65931), .Q(n38550) );
  IMUX40 U44014 ( .A(n65656), .B(\OFill[29][0] ), .C(n65658), .D(n65659), .S0(
        n65821), .S1(n65931), .Q(n38553) );
  IMUX40 U44015 ( .A(n65652), .B(\OFill[25][0] ), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65813), .S1(n65931), .Q(n38551) );
  IMUX40 U43848 ( .A(n38550), .B(n38551), .C(n38552), .D(n38553), .S0(N1018), 
        .S1(N1017), .Q(n38549) );
  IMUX40 U46705 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65785), .S1(n65926), .Q(n41110) );
  IMUX40 U46702 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65809), .S1(n65926), .Q(n41113) );
  IMUX40 U46703 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65793), .S1(n65926), .Q(n41111) );
  IMUX40 U46536 ( .A(n41110), .B(n41111), .C(n41112), .D(n41113), .S0(N1042), 
        .S1(N1041), .Q(n41109) );
  IMUX40 U46033 ( .A(n65644), .B(\OFill[17][0] ), .C(n65646), .D(n65647), .S0(
        n65792), .S1(n65928), .Q(n40470) );
  IMUX40 U46030 ( .A(n65656), .B(\OFill[29][0] ), .C(\OFill[30][0] ), .D(
        n65659), .S0(n65793), .S1(n65928), .Q(n40473) );
  IMUX40 U46031 ( .A(n65652), .B(n65653), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65793), .S1(n65928), .Q(n40471) );
  IMUX40 U45864 ( .A(n40470), .B(n40471), .C(n40472), .D(n40473), .S0(N1036), 
        .S1(N1035), .Q(n40469) );
  IMUX40 U47377 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65797), .S1(n65924), .Q(n41750) );
  IMUX40 U47374 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65797), .S1(n65924), .Q(n41753) );
  IMUX40 U47375 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65797), .S1(n65924), .Q(n41751) );
  IMUX40 U47208 ( .A(n41750), .B(n41751), .C(n41752), .D(n41753), .S0(N1048), 
        .S1(N1047), .Q(n41749) );
  IMUX40 U48725 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65829), .S1(N1082), .Q(n43035) );
  IMUX40 U48722 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65824), .S1(N1082), .Q(n43038) );
  IMUX40 U48723 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65825), .S1(n65923), .Q(n43036) );
  IMUX40 U48553 ( .A(n43035), .B(n43036), .C(n43037), .D(n43038), .S0(N1060), 
        .S1(N1059), .Q(n43034) );
  IMUX40 U48721 ( .A(\OFill[16][0] ), .B(n65645), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65786), .S1(n65922), .Q(n43030) );
  IMUX40 U48718 ( .A(\OFill[28][0] ), .B(n65657), .C(\OFill[30][0] ), .D(
        \OFill[31][0] ), .S0(n65822), .S1(n65911), .Q(n43033) );
  IMUX40 U48719 ( .A(\OFill[24][0] ), .B(n65653), .C(n65654), .D(n65655), .S0(
        n65823), .S1(n65923), .Q(n43031) );
  IMUX40 U48552 ( .A(n43030), .B(n43031), .C(n43032), .D(n43033), .S0(N1060), 
        .S1(N1059), .Q(n43029) );
  IMUX40 U48053 ( .A(n65660), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65833), .S1(n65781), .Q(n42395) );
  IMUX40 U48050 ( .A(n65672), .B(n65673), .C(\OFill[14][0] ), .D(
        \OFill[15][0] ), .S0(n65832), .S1(n65778), .Q(n42398) );
  IMUX40 U48051 ( .A(n65668), .B(\OFill[9][0] ), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65832), .S1(n65781), .Q(n42396) );
  IMUX40 U47881 ( .A(n42395), .B(n42396), .C(n42397), .D(n42398), .S0(N1054), 
        .S1(N1053), .Q(n42394) );
  IMUX40 U48049 ( .A(n65644), .B(n65645), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65832), .S1(n65775), .Q(n42390) );
  IMUX40 U48046 ( .A(n65656), .B(n65657), .C(\OFill[30][0] ), .D(
        \OFill[31][0] ), .S0(n65848), .S1(n65780), .Q(n42393) );
  IMUX40 U48047 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65899), 
        .S1(n65767), .Q(n42391) );
  IMUX40 U47880 ( .A(n42390), .B(n42391), .C(n42392), .D(n42393), .S0(N1054), 
        .S1(N1053), .Q(n42389) );
  IMUX40 U49393 ( .A(n65644), .B(\OFill[17][0] ), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65907), .S1(n65749), .Q(n43670) );
  IMUX40 U49390 ( .A(n65656), .B(\OFill[29][0] ), .C(\OFill[30][0] ), .D(
        \OFill[31][0] ), .S0(n65904), .S1(N1208), .Q(n43673) );
  IMUX40 U49391 ( .A(n65652), .B(\OFill[25][0] ), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65880), .S1(n65752), .Q(n43671) );
  IMUX40 U49224 ( .A(n43670), .B(n43671), .C(n43672), .D(n43673), .S0(N1066), 
        .S1(n65920), .Q(n43669) );
  IMUX40 U50741 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65880), .S1(n65774), .Q(n44955) );
  IMUX40 U50738 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65857), .S1(n65775), .Q(n44958) );
  IMUX40 U50739 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65854), .S1(n65768), .Q(n44956) );
  IMUX40 U50569 ( .A(n44955), .B(n44956), .C(n44957), .D(n44958), .S0(N1078), 
        .S1(N1077), .Q(n44954) );
  IMUX40 U50737 ( .A(\OFill[16][0] ), .B(n65645), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65833), .S1(n65777), .Q(n44950) );
  IMUX40 U50734 ( .A(\OFill[28][0] ), .B(n65657), .C(\OFill[30][0] ), .D(
        \OFill[31][0] ), .S0(n65887), .S1(n65774), .Q(n44953) );
  IMUX40 U50735 ( .A(\OFill[24][0] ), .B(n65653), .C(n65654), .D(n65655), .S0(
        n65901), .S1(n65761), .Q(n44951) );
  IMUX40 U50568 ( .A(n44950), .B(n44951), .C(n44952), .D(n44953), .S0(N1078), 
        .S1(N1077), .Q(n44949) );
  IMUX40 U51409 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65821), .S1(n65922), .Q(n45590) );
  IMUX40 U51406 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65820), .S1(n65922), .Q(n45593) );
  IMUX40 U51407 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65820), .S1(n65922), .Q(n45591) );
  IMUX40 U51240 ( .A(n45590), .B(n45591), .C(n45592), .D(n45593), .S0(N1084), 
        .S1(N1083), .Q(n45589) );
  IMUX40 U64853 ( .A(\OFill[0][0] ), .B(n65661), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65794), .S1(n65911), .Q(n58395) );
  IMUX40 U64850 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(n65674), .D(
        \OFill[15][0] ), .S0(n65796), .S1(n65911), .Q(n58398) );
  IMUX40 U64851 ( .A(\OFill[8][0] ), .B(n65669), .C(\OFill[10][0] ), .D(
        \OFill[11][0] ), .S0(n65797), .S1(n65911), .Q(n58396) );
  IMUX40 U64681 ( .A(n58395), .B(n58396), .C(n58397), .D(n58398), .S0(N1204), 
        .S1(N1203), .Q(n58394) );
  IMUX40 U64849 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(n65646), .D(
        n65647), .S0(n65792), .S1(n65911), .Q(n58390) );
  IMUX40 U64846 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(n65659), .S0(n65822), .S1(n65911), .Q(n58393) );
  IMUX40 U64847 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65791), .S1(n65911), .Q(n58391) );
  IMUX40 U64680 ( .A(n58390), .B(n58391), .C(n58392), .D(n58393), .S0(N1204), 
        .S1(N1203), .Q(n58389) );
  IMUX40 U64177 ( .A(n65644), .B(\OFill[17][0] ), .C(n65646), .D(n65647), .S0(
        n65903), .S1(n65771), .Q(n57750) );
  IMUX40 U64174 ( .A(n65656), .B(\OFill[29][0] ), .C(\OFill[30][0] ), .D(
        n65659), .S0(n65893), .S1(n65769), .Q(n57753) );
  IMUX40 U64175 ( .A(n65652), .B(\OFill[25][0] ), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65857), .S1(n65765), .Q(n57751) );
  IMUX40 U64008 ( .A(n57750), .B(n57751), .C(n57752), .D(n57753), .S0(N1198), 
        .S1(N1197), .Q(n57749) );
  IMUX40 U65521 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65888), .S1(n65755), .Q(n59030) );
  IMUX40 U65518 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65890), .S1(n65750), .Q(n59033) );
  IMUX40 U65519 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65893), .S1(n65757), .Q(n59031) );
  IMUX40 U65352 ( .A(n59030), .B(n59031), .C(n59032), .D(n59033), .S0(N1210), 
        .S1(n65919), .Q(n59029) );
  IMUX40 U15797 ( .A(n65724), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65859), .S1(n65768), .Q(n11675) );
  IMUX40 U15794 ( .A(n65736), .B(\GFill[13][0] ), .C(\GFill[14][0] ), .D(
        \GFill[15][0] ), .S0(n65860), .S1(n65780), .Q(n11678) );
  IMUX40 U15795 ( .A(n65732), .B(\GFill[9][0] ), .C(\GFill[10][0] ), .D(
        \GFill[11][0] ), .S0(n65859), .S1(n65779), .Q(n11676) );
  IMUX40 U15625 ( .A(n11675), .B(n11676), .C(n11677), .D(n11678), .S0(N1054), 
        .S1(N1053), .Q(n11674) );
  IMUX40 U15793 ( .A(n65708), .B(n65709), .C(n65710), .D(\GFill[19][0] ), .S0(
        n65860), .S1(n65779), .Q(n11670) );
  IMUX40 U15790 ( .A(n65720), .B(n65721), .C(n65722), .D(\GFill[31][0] ), .S0(
        n65861), .S1(n65775), .Q(n11673) );
  IMUX40 U15791 ( .A(n65716), .B(n65717), .C(n65718), .D(\GFill[27][0] ), .S0(
        n65861), .S1(n65781), .Q(n11671) );
  IMUX40 U15624 ( .A(n11670), .B(n11671), .C(n11672), .D(n11673), .S0(N1054), 
        .S1(N1053), .Q(n11669) );
  IMUX40 U17137 ( .A(\GFill[16][0] ), .B(n65709), .C(n65710), .D(
        \GFill[19][0] ), .S0(n65858), .S1(n65755), .Q(n12950) );
  IMUX40 U17134 ( .A(\GFill[28][0] ), .B(n65721), .C(n65722), .D(
        \GFill[31][0] ), .S0(n65857), .S1(n65752), .Q(n12953) );
  IMUX40 U17135 ( .A(\GFill[24][0] ), .B(n65717), .C(n65718), .D(
        \GFill[27][0] ), .S0(n65857), .S1(n65745), .Q(n12951) );
  IMUX40 U16968 ( .A(n12950), .B(n12951), .C(n12952), .D(n12953), .S0(N1066), 
        .S1(n65920), .Q(n12949) );
  IMUX40 U16465 ( .A(n65708), .B(\GFill[17][0] ), .C(\GFill[18][0] ), .D(
        \GFill[19][0] ), .S0(n65812), .S1(n65922), .Q(n12310) );
  IMUX40 U16462 ( .A(n65720), .B(\GFill[29][0] ), .C(\GFill[30][0] ), .D(
        \GFill[31][0] ), .S0(n65786), .S1(n65912), .Q(n12313) );
  IMUX40 U16463 ( .A(n65716), .B(\GFill[25][0] ), .C(\GFill[26][0] ), .D(
        \GFill[27][0] ), .S0(n65802), .S1(n65537), .Q(n12311) );
  IMUX40 U16296 ( .A(n12310), .B(n12311), .C(n12312), .D(n12313), .S0(N1060), 
        .S1(N1059), .Q(n12309) );
  IMUX40 U18481 ( .A(\GFill[16][0] ), .B(n65709), .C(n65710), .D(
        \GFill[19][0] ), .S0(n65907), .S1(n65773), .Q(n14230) );
  IMUX40 U18478 ( .A(\GFill[28][0] ), .B(n65721), .C(n65722), .D(
        \GFill[31][0] ), .S0(n65877), .S1(n65771), .Q(n14233) );
  IMUX40 U18479 ( .A(\GFill[24][0] ), .B(n65717), .C(n65718), .D(
        \GFill[27][0] ), .S0(n65851), .S1(n65777), .Q(n14231) );
  IMUX40 U18312 ( .A(n14230), .B(n14231), .C(n14232), .D(n14233), .S0(N1078), 
        .S1(N1077), .Q(n14229) );
  IMUX40 U19153 ( .A(n65708), .B(\GFill[17][0] ), .C(\GFill[18][0] ), .D(
        \GFill[19][0] ), .S0(n65807), .S1(n65923), .Q(n14870) );
  IMUX40 U19150 ( .A(n65720), .B(\GFill[29][0] ), .C(\GFill[30][0] ), .D(
        \GFill[31][0] ), .S0(n65816), .S1(N1082), .Q(n14873) );
  IMUX40 U19151 ( .A(n65716), .B(\GFill[25][0] ), .C(\GFill[26][0] ), .D(
        \GFill[27][0] ), .S0(n65806), .S1(n65912), .Q(n14871) );
  IMUX40 U18984 ( .A(n14870), .B(n14871), .C(n14872), .D(n14873), .S0(N1084), 
        .S1(N1083), .Q(n14869) );
  IMUX40 U32593 ( .A(n65708), .B(\GFill[17][0] ), .C(\GFill[18][0] ), .D(
        n65711), .S0(n65831), .S1(n65911), .Q(n27670) );
  IMUX40 U32590 ( .A(n65720), .B(\GFill[29][0] ), .C(\GFill[30][0] ), .D(
        n65723), .S0(n65806), .S1(n65743), .Q(n27673) );
  IMUX40 U32591 ( .A(n65716), .B(\GFill[25][0] ), .C(\GFill[26][0] ), .D(
        n65719), .S0(n65827), .S1(N1082), .Q(n27671) );
  IMUX40 U32424 ( .A(n27670), .B(n27671), .C(n27672), .D(n27673), .S0(N1204), 
        .S1(N1203), .Q(n27669) );
  IMUX40 U31921 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(n65711), .S0(n65903), .S1(n65779), .Q(n27030) );
  IMUX40 U31918 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(n65723), .S0(n65836), .S1(n65760), .Q(n27033) );
  IMUX40 U31919 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(n65719), .S0(n65855), .S1(n65780), .Q(n27031) );
  IMUX40 U31752 ( .A(n27030), .B(n27031), .C(n27032), .D(n27033), .S0(N1198), 
        .S1(N1197), .Q(n27029) );
  IMUX40 U33265 ( .A(n65708), .B(\GFill[17][0] ), .C(\GFill[18][0] ), .D(
        \GFill[19][0] ), .S0(n65884), .S1(n65744), .Q(n28310) );
  IMUX40 U33262 ( .A(n65720), .B(\GFill[29][0] ), .C(\GFill[30][0] ), .D(
        \GFill[31][0] ), .S0(n65837), .S1(n65745), .Q(n28313) );
  IMUX40 U33263 ( .A(n65716), .B(\GFill[25][0] ), .C(\GFill[26][0] ), .D(
        \GFill[27][0] ), .S0(n65896), .S1(n65744), .Q(n28311) );
  IMUX40 U33096 ( .A(n28310), .B(n28311), .C(n28312), .D(n28313), .S0(N1210), 
        .S1(n65919), .Q(n28309) );
  IMUX40 U34613 ( .A(\GFill[0][0] ), .B(n65725), .C(n65726), .D(n65727), .S0(
        n65782), .S1(n65911), .Q(n29595) );
  IMUX40 U34610 ( .A(\GFill[12][0] ), .B(n65737), .C(n65738), .D(n65739), .S0(
        n65808), .S1(N1130), .Q(n29598) );
  IMUX40 U34611 ( .A(\GFill[8][0] ), .B(n65733), .C(n65734), .D(n65735), .S0(
        n65808), .S1(N1148), .Q(n29596) );
  IMUX40 U34441 ( .A(n29595), .B(n29596), .C(n29597), .D(n29598), .S0(N1222), 
        .S1(N1221), .Q(n29594) );
  IMUX40 U34609 ( .A(\GFill[16][0] ), .B(n65709), .C(n65710), .D(n65711), .S0(
        n65808), .S1(N1220), .Q(n29590) );
  IMUX40 U34606 ( .A(\GFill[28][0] ), .B(n65721), .C(n65722), .D(n65723), .S0(
        n65808), .S1(n65538), .Q(n29593) );
  IMUX40 U34607 ( .A(\GFill[24][0] ), .B(n65717), .C(n65718), .D(n65719), .S0(
        n65808), .S1(N1148), .Q(n29591) );
  IMUX40 U34440 ( .A(n29590), .B(n29591), .C(n29592), .D(n29593), .S0(N1222), 
        .S1(N1221), .Q(n29589) );
  IMUX40 U33941 ( .A(\GFill[0][0] ), .B(n65725), .C(n65726), .D(n65727), .S0(
        n65903), .S1(n65780), .Q(n28955) );
  IMUX40 U33938 ( .A(\GFill[12][0] ), .B(n65737), .C(n65738), .D(n65739), .S0(
        n65897), .S1(n65760), .Q(n28958) );
  IMUX40 U33939 ( .A(\GFill[8][0] ), .B(n65733), .C(n65734), .D(n65735), .S0(
        n65877), .S1(n65776), .Q(n28956) );
  IMUX40 U33769 ( .A(n28955), .B(n28956), .C(n28957), .D(n28958), .S0(N1216), 
        .S1(N1215), .Q(n28954) );
  IMUX40 U33937 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65840), 
        .S1(n65760), .Q(n28950) );
  IMUX40 U33934 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65873), 
        .S1(n65760), .Q(n28953) );
  IMUX40 U33935 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65846), 
        .S1(n65760), .Q(n28951) );
  IMUX40 U33768 ( .A(n28950), .B(n28951), .C(n28952), .D(n28953), .S0(N1216), 
        .S1(N1215), .Q(n28949) );
  IMUX40 U66869 ( .A(\OFill[0][0] ), .B(n65661), .C(n65662), .D(n65663), .S0(
        n65785), .S1(n65743), .Q(n60315) );
  IMUX40 U66866 ( .A(n65672), .B(n65673), .C(n65674), .D(n65675), .S0(n65813), 
        .S1(n65743), .Q(n60318) );
  IMUX40 U66867 ( .A(n65668), .B(n65669), .C(n65670), .D(n65671), .S0(n65815), 
        .S1(n65743), .Q(n60316) );
  IMUX40 U66697 ( .A(n60315), .B(n60316), .C(n60317), .D(n60318), .S0(N1222), 
        .S1(N1221), .Q(n60314) );
  IMUX40 U66865 ( .A(\OFill[16][0] ), .B(n65645), .C(n65646), .D(n65647), .S0(
        n65810), .S1(n65743), .Q(n60310) );
  IMUX40 U66862 ( .A(\OFill[28][0] ), .B(n65657), .C(n65658), .D(n65659), .S0(
        n65812), .S1(n65743), .Q(n60313) );
  IMUX40 U66863 ( .A(\OFill[24][0] ), .B(n65653), .C(n65654), .D(n65655), .S0(
        n65799), .S1(n65743), .Q(n60311) );
  IMUX40 U66696 ( .A(n60310), .B(n60311), .C(n60312), .D(n60313), .S0(N1222), 
        .S1(N1221), .Q(n60309) );
  IMUX40 U66197 ( .A(\OFill[0][0] ), .B(n65661), .C(n65662), .D(n65663), .S0(
        n65844), .S1(n65764), .Q(n59675) );
  IMUX40 U66194 ( .A(\OFill[12][0] ), .B(n65673), .C(n65674), .D(n65675), .S0(
        n65908), .S1(n65764), .Q(n59678) );
  IMUX40 U66195 ( .A(\OFill[8][0] ), .B(n65669), .C(n65670), .D(n65671), .S0(
        n65869), .S1(n65764), .Q(n59676) );
  IMUX40 U66025 ( .A(n59675), .B(n59676), .C(n59677), .D(n59678), .S0(N1216), 
        .S1(N1215), .Q(n59674) );
  IMUX40 U66193 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65846), 
        .S1(n65764), .Q(n59670) );
  IMUX40 U66190 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65898), 
        .S1(n65763), .Q(n59673) );
  IMUX40 U66191 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(N1207), 
        .S1(n65763), .Q(n59671) );
  IMUX40 U66024 ( .A(n59670), .B(n59671), .C(n59672), .D(n59673), .S0(N1216), 
        .S1(N1215), .Q(n59669) );
  IMUX40 U35953 ( .A(n65708), .B(n65709), .C(n65710), .D(n65711), .S0(n65886), 
        .S1(n65776), .Q(n30870) );
  IMUX40 U35950 ( .A(n65720), .B(n65721), .C(n65722), .D(n65723), .S0(n65860), 
        .S1(n65765), .Q(n30873) );
  IMUX40 U35951 ( .A(n65716), .B(n65717), .C(n65718), .D(n65719), .S0(n65861), 
        .S1(n65760), .Q(n30871) );
  IMUX40 U35784 ( .A(n30870), .B(n30871), .C(n30872), .D(n30873), .S0(N1234), 
        .S1(N1233), .Q(n30869) );
  IMUX40 U68209 ( .A(n65644), .B(n65645), .C(n65646), .D(n65647), .S0(n65904), 
        .S1(n65764), .Q(n61590) );
  IMUX40 U68206 ( .A(n65656), .B(n65657), .C(n65658), .D(n65659), .S0(n65865), 
        .S1(n65763), .Q(n61593) );
  IMUX40 U68207 ( .A(n65652), .B(n65653), .C(n65654), .D(n65655), .S0(n65900), 
        .S1(n65759), .Q(n61591) );
  IMUX40 U68040 ( .A(n61590), .B(n61591), .C(n61592), .D(n61593), .S0(N1234), 
        .S1(N1233), .Q(n61589) );
  IMUX40 U63505 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(n65646), .D(
        n65647), .S0(n65832), .S1(n65760), .Q(n57110) );
  IMUX40 U63502 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(n65659), .S0(n65899), .S1(n65765), .Q(n57113) );
  IMUX40 U63503 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(n65655), .S0(n65832), .S1(n65763), .Q(n57111) );
  IMUX40 U63336 ( .A(n57110), .B(n57111), .C(n57112), .D(n57113), .S0(N1192), 
        .S1(N1191), .Q(n57109) );
  IMUX40 U31249 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(n65711), .S0(n65873), .S1(n65772), .Q(n26390) );
  IMUX40 U31246 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(n65723), .S0(n65868), .S1(n65781), .Q(n26393) );
  IMUX40 U31247 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(n65719), .S0(n65901), .S1(n65779), .Q(n26391) );
  IMUX40 U31080 ( .A(n26390), .B(n26391), .C(n26392), .D(n26393), .S0(N1192), 
        .S1(N1191), .Q(n26389) );
  IMUX40 U21845 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65844), .S1(n65780), .Q(n17435) );
  IMUX40 U21842 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65845), .S1(n65764), .Q(n17438) );
  IMUX40 U21843 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65845), .S1(n65763), .Q(n17436) );
  IMUX40 U21673 ( .A(n17435), .B(n17436), .C(n17437), .D(n17438), .S0(N1108), 
        .S1(N1107), .Q(n17434) );
  IMUX40 U21841 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65845), .S1(n65765), .Q(n17430) );
  IMUX40 U21838 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65846), .S1(n65760), .Q(n17433) );
  IMUX40 U21839 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65846), .S1(n65781), .Q(n17431) );
  IMUX40 U21672 ( .A(n17430), .B(n17431), .C(n17432), .D(n17433), .S0(N1108), 
        .S1(N1107), .Q(n17429) );
  IMUX40 U54097 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65853), .S1(n65775), .Q(n48150) );
  IMUX40 U54094 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65852), .S1(n65769), .Q(n48153) );
  IMUX40 U54095 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65853), .S1(n65761), .Q(n48151) );
  IMUX40 U53928 ( .A(n48150), .B(n48151), .C(n48152), .D(n48153), .S0(N1108), 
        .S1(N1107), .Q(n48149) );
  IMUX40 U50065 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65842), .S1(n65756), .Q(n44310) );
  IMUX40 U50062 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65841), .S1(n65755), .Q(n44313) );
  IMUX40 U50063 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65842), .S1(n65745), .Q(n44311) );
  IMUX40 U49896 ( .A(n44310), .B(n44311), .C(n44312), .D(n44313), .S0(N1072), 
        .S1(n65918), .Q(n44309) );
  IMUX40 U62161 ( .A(n65644), .B(\OFill[17][0] ), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65868), .S1(n65748), .Q(n55830) );
  IMUX40 U62158 ( .A(n65656), .B(\OFill[29][0] ), .C(\OFill[30][0] ), .D(
        \OFill[31][0] ), .S0(n65867), .S1(n65747), .Q(n55833) );
  IMUX40 U62159 ( .A(n65652), .B(\OFill[25][0] ), .C(\OFill[26][0] ), .D(
        \OFill[27][0] ), .S0(n65868), .S1(n65750), .Q(n55831) );
  IMUX40 U61992 ( .A(n55830), .B(n55831), .C(n55832), .D(n55833), .S0(N1180), 
        .S1(n65915), .Q(n55829) );
  IMUX40 U17809 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65835), .S1(n65747), .Q(n13590) );
  IMUX40 U17806 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65836), .S1(n65750), .Q(n13593) );
  IMUX40 U17807 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65835), .S1(n65756), .Q(n13591) );
  IMUX40 U17640 ( .A(n13590), .B(n13591), .C(n13592), .D(n13593), .S0(N1072), 
        .S1(n65918), .Q(n13589) );
  IMUX40 U29905 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65904), .S1(n65745), .Q(n25110) );
  IMUX40 U29902 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65853), .S1(n65752), .Q(n25113) );
  IMUX40 U29903 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65877), .S1(n65752), .Q(n25111) );
  IMUX40 U29736 ( .A(n25110), .B(n25111), .C(n25112), .D(n25113), .S0(N1180), 
        .S1(n65916), .Q(n25109) );
  IMUX40 U28565 ( .A(\GFill[0][0] ), .B(\GFill[1][0] ), .C(\GFill[2][0] ), .D(
        \GFill[3][0] ), .S0(n65881), .S1(n65757), .Q(n23835) );
  IMUX40 U28562 ( .A(\GFill[12][0] ), .B(\GFill[13][0] ), .C(\GFill[14][0] ), 
        .D(\GFill[15][0] ), .S0(n65870), .S1(n65751), .Q(n23838) );
  IMUX40 U28563 ( .A(\GFill[8][0] ), .B(\GFill[9][0] ), .C(\GFill[10][0] ), 
        .D(\GFill[11][0] ), .S0(n65870), .S1(n65751), .Q(n23836) );
  IMUX40 U28393 ( .A(n23835), .B(n23836), .C(n23837), .D(n23838), .S0(N1168), 
        .S1(n65915), .Q(n23834) );
  IMUX40 U28561 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(n65710), .D(
        \GFill[19][0] ), .S0(n65870), .S1(n65751), .Q(n23830) );
  IMUX40 U28558 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(n65722), .D(
        \GFill[31][0] ), .S0(n65871), .S1(n65751), .Q(n23833) );
  IMUX40 U28559 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(n65718), .D(
        \GFill[27][0] ), .S0(n65871), .S1(n65751), .Q(n23831) );
  IMUX40 U28392 ( .A(n23830), .B(n23831), .C(n23832), .D(n23833), .S0(N1168), 
        .S1(n65916), .Q(n23829) );
  IMUX40 U27217 ( .A(\GFill[16][0] ), .B(\GFill[17][0] ), .C(\GFill[18][0] ), 
        .D(\GFill[19][0] ), .S0(n65842), .S1(n65746), .Q(n22550) );
  IMUX40 U27214 ( .A(\GFill[28][0] ), .B(\GFill[29][0] ), .C(\GFill[30][0] ), 
        .D(\GFill[31][0] ), .S0(n65885), .S1(n65746), .Q(n22553) );
  IMUX40 U27215 ( .A(\GFill[24][0] ), .B(\GFill[25][0] ), .C(\GFill[26][0] ), 
        .D(\GFill[27][0] ), .S0(n65889), .S1(n65746), .Q(n22551) );
  IMUX40 U27048 ( .A(n22550), .B(n22551), .C(n22552), .D(n22553), .S0(N1156), 
        .S1(n65917), .Q(n22549) );
  IMUX40 U60821 ( .A(\OFill[0][0] ), .B(\OFill[1][0] ), .C(\OFill[2][0] ), .D(
        \OFill[3][0] ), .S0(n65847), .S1(n65749), .Q(n54555) );
  IMUX40 U60818 ( .A(\OFill[12][0] ), .B(\OFill[13][0] ), .C(\OFill[14][0] ), 
        .D(\OFill[15][0] ), .S0(n65910), .S1(n65750), .Q(n54558) );
  IMUX40 U60819 ( .A(\OFill[8][0] ), .B(\OFill[9][0] ), .C(\OFill[10][0] ), 
        .D(\OFill[11][0] ), .S0(n65849), .S1(n65749), .Q(n54556) );
  IMUX40 U60649 ( .A(n54555), .B(n54556), .C(n54557), .D(n54558), .S0(N1168), 
        .S1(n65917), .Q(n54554) );
  IMUX40 U60817 ( .A(\OFill[16][0] ), .B(n65645), .C(\OFill[18][0] ), .D(
        \OFill[19][0] ), .S0(n65853), .S1(n65750), .Q(n54550) );
  IMUX40 U60814 ( .A(\OFill[28][0] ), .B(n65657), .C(n65658), .D(
        \OFill[31][0] ), .S0(n65909), .S1(n65750), .Q(n54553) );
  IMUX40 U60815 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(n65654), .D(
        n65655), .S0(n65854), .S1(n65750), .Q(n54551) );
  IMUX40 U60648 ( .A(n54550), .B(n54551), .C(n54552), .D(n54553), .S0(N1168), 
        .S1(n65916), .Q(n54549) );
  IMUX40 U59473 ( .A(\OFill[16][0] ), .B(\OFill[17][0] ), .C(\OFill[18][0] ), 
        .D(\OFill[19][0] ), .S0(n65875), .S1(n65744), .Q(n53270) );
  IMUX40 U59470 ( .A(\OFill[28][0] ), .B(\OFill[29][0] ), .C(\OFill[30][0] ), 
        .D(\OFill[31][0] ), .S0(n65837), .S1(n65745), .Q(n53273) );
  IMUX40 U59471 ( .A(\OFill[24][0] ), .B(\OFill[25][0] ), .C(\OFill[26][0] ), 
        .D(\OFill[27][0] ), .S0(n65866), .S1(n65744), .Q(n53271) );
  IMUX40 U59304 ( .A(n53270), .B(n53271), .C(n53272), .D(n53273), .S0(N1156), 
        .S1(n65918), .Q(n53269) );
  MUX41 U28394 ( .A(n23834), .B(n23824), .C(n23829), .D(n23819), .S0(N1170), 
        .S1(N1169), .Q(N4400) );
  MUX41 U60650 ( .A(n54554), .B(n54544), .C(n54549), .D(n54539), .S0(N1170), 
        .S1(N1169), .Q(N6670) );
  IMUX40 U23017 ( .A(n18715), .B(n18716), .C(n18717), .D(n18718), .S0(N1120), 
        .S1(n65917), .Q(n18714) );
  IMUX40 U23014 ( .A(n18700), .B(n18701), .C(n18702), .D(n18703), .S0(N11412), 
        .S1(n65917), .Q(n18699) );
  IMUX40 U23015 ( .A(n18705), .B(n18706), .C(n18707), .D(n18708), .S0(N1120), 
        .S1(n65917), .Q(n18704) );
  MUX41 U23018 ( .A(n18714), .B(n18704), .C(n18709), .D(n18699), .S0(N1122), 
        .S1(N1121), .Q(N4020) );
  IMUX40 U70729 ( .A(n64155), .B(n64156), .C(n64157), .D(n64158), .S0(N1258), 
        .S1(N1257), .Q(n64154) );
  IMUX40 U70726 ( .A(n64140), .B(n64141), .C(n64142), .D(n64143), .S0(N1258), 
        .S1(N1257), .Q(n64139) );
  IMUX40 U70727 ( .A(n64145), .B(n64146), .C(n64147), .D(n64148), .S0(N1258), 
        .S1(N1257), .Q(n64144) );
  MUX41 U70730 ( .A(n64154), .B(n64144), .C(n64149), .D(n64139), .S0(N1260), 
        .S1(N1259), .Q(N7360) );
  IMUX40 U8902 ( .A(n5260), .B(n5261), .C(n5262), .D(n5263), .S0(N706), .S1(
        N705), .Q(n5259) );
  IMUX40 U8903 ( .A(n5265), .B(n5266), .C(n5267), .D(n5268), .S0(N706), .S1(
        N705), .Q(n5264) );
  MUX41 U8906 ( .A(n5274), .B(n5264), .C(n5269), .D(n5259), .S0(N708), .S1(
        N707), .Q(N3040) );
  IMUX40 U42502 ( .A(n37260), .B(n37261), .C(n37262), .D(n37263), .S0(N1006), 
        .S1(N1005), .Q(n37259) );
  IMUX40 U42503 ( .A(n37265), .B(n37266), .C(n37267), .D(n37268), .S0(N1006), 
        .S1(N1005), .Q(n37264) );
  MUX41 U42506 ( .A(n37274), .B(n37264), .C(n37269), .D(n37259), .S0(N1008), 
        .S1(N1007), .Q(N5432) );
  IMUX40 U62665 ( .A(n56475), .B(n56476), .C(n56477), .D(n56478), .S0(N1186), 
        .S1(N1185), .Q(n56474) );
  IMUX40 U62662 ( .A(n56460), .B(n56461), .C(n56462), .D(n56463), .S0(N1186), 
        .S1(N1185), .Q(n56459) );
  IMUX40 U62663 ( .A(n56465), .B(n56466), .C(n56467), .D(n56468), .S0(N1186), 
        .S1(N1185), .Q(n56464) );
  MUX41 U62666 ( .A(n56474), .B(n56464), .C(n56469), .D(n56459), .S0(N1188), 
        .S1(N1187), .Q(N6809) );
  IMUX40 U16969 ( .A(n12955), .B(n12956), .C(n12957), .D(n12958), .S0(N1066), 
        .S1(n65919), .Q(n12954) );
  IMUX40 U16966 ( .A(n12940), .B(n12941), .C(n12942), .D(n12943), .S0(N1066), 
        .S1(n65920), .Q(n12939) );
  IMUX40 U16967 ( .A(n12945), .B(n12946), .C(n12947), .D(n12948), .S0(N1066), 
        .S1(n65919), .Q(n12944) );
  MUX41 U16970 ( .A(n12954), .B(n12944), .C(n12949), .D(n12939), .S0(N1068), 
        .S1(N1067), .Q(N3631) );
  IMUX40 U14953 ( .A(n11035), .B(n11036), .C(n11037), .D(n11038), .S0(N1048), 
        .S1(N1047), .Q(n11034) );
  IMUX40 U14950 ( .A(n11020), .B(n11021), .C(n11022), .D(n11023), .S0(N1048), 
        .S1(N1047), .Q(n11019) );
  IMUX40 U14951 ( .A(n11025), .B(n11026), .C(n11027), .D(n11028), .S0(N1048), 
        .S1(N1047), .Q(n11024) );
  MUX41 U14954 ( .A(n11034), .B(n11024), .C(n11029), .D(n11019), .S0(N1050), 
        .S1(N1049), .Q(N3504) );
  IMUX40 U44521 ( .A(n39195), .B(n39196), .C(n39197), .D(n39198), .S0(N1024), 
        .S1(N1023), .Q(n39194) );
  IMUX40 U44518 ( .A(n39180), .B(n39181), .C(n39182), .D(n39183), .S0(N1024), 
        .S1(N1023), .Q(n39179) );
  IMUX40 U44519 ( .A(n39185), .B(n39186), .C(n39187), .D(n39188), .S0(N1024), 
        .S1(N1023), .Q(n39184) );
  MUX41 U44522 ( .A(n39194), .B(n39184), .C(n39189), .D(n39179), .S0(N1026), 
        .S1(N1025), .Q(N5587) );
  IMUX40 U46537 ( .A(n41115), .B(n41116), .C(n41117), .D(n41118), .S0(N1042), 
        .S1(N1041), .Q(n41114) );
  IMUX40 U46534 ( .A(n41100), .B(n41101), .C(n41102), .D(n41103), .S0(N1042), 
        .S1(N1041), .Q(n41099) );
  IMUX40 U46535 ( .A(n41105), .B(n41106), .C(n41107), .D(n41108), .S0(N1042), 
        .S1(N1041), .Q(n41104) );
  MUX41 U46538 ( .A(n41114), .B(n41104), .C(n41109), .D(n41099), .S0(N1044), 
        .S1(N1043), .Q(N5742) );
  IMUX40 U8233 ( .A(n4635), .B(n4636), .C(n4637), .D(n4638), .S0(N700), .S1(
        N699), .Q(n4634) );
  IMUX40 U8230 ( .A(n4620), .B(n4621), .C(n4622), .D(n4623), .S0(N700), .S1(
        N699), .Q(n4619) );
  IMUX40 U8231 ( .A(n4625), .B(n4626), .C(n4627), .D(n4628), .S0(N700), .S1(
        N699), .Q(n4624) );
  MUX41 U8234 ( .A(n4634), .B(n4624), .C(n4629), .D(n4619), .S0(N702), .S1(
        N701), .Q(N3008) );
  IMUX40 U10918 ( .A(n7180), .B(n7181), .C(n7182), .D(n7183), .S0(N724), .S1(
        N723), .Q(n7179) );
  IMUX40 U10919 ( .A(n7185), .B(n7186), .C(n7187), .D(n7188), .S0(N724), .S1(
        N723), .Q(n7184) );
  MUX41 U10922 ( .A(n7194), .B(n7184), .C(n7189), .D(n7179), .S0(N726), .S1(
        N725), .Q(N3194) );
  IMUX40 U27718 ( .A(n23180), .B(n23181), .C(n23182), .D(n23183), .S0(N874), 
        .S1(N873), .Q(n23179) );
  IMUX40 U27719 ( .A(n23185), .B(n23186), .C(n23187), .D(n23188), .S0(N874), 
        .S1(N873), .Q(n23184) );
  MUX41 U27722 ( .A(n23194), .B(n23184), .C(n23189), .D(n23179), .S0(N876), 
        .S1(N875), .Q(N4368) );
  IMUX40 U25702 ( .A(n21260), .B(n21261), .C(n21262), .D(n21263), .S0(N856), 
        .S1(N855), .Q(n21259) );
  IMUX40 U25703 ( .A(n21265), .B(n21266), .C(n21267), .D(n21268), .S0(N856), 
        .S1(N855), .Q(n21264) );
  MUX41 U25706 ( .A(n21274), .B(n21264), .C(n21269), .D(n21259), .S0(N858), 
        .S1(N857), .Q(N4229) );
  IMUX40 U59974 ( .A(n53900), .B(n53901), .C(n53902), .D(n53903), .S0(N1162), 
        .S1(N1161), .Q(n53899) );
  IMUX40 U59975 ( .A(n53905), .B(n53906), .C(n53907), .D(n53908), .S0(N1162), 
        .S1(N1161), .Q(n53904) );
  MUX41 U59978 ( .A(n53914), .B(n53904), .C(n53909), .D(n53899), .S0(N1164), 
        .S1(N1163), .Q(N6638) );
  IMUX40 U57958 ( .A(n51980), .B(n51981), .C(n51982), .D(n51983), .S0(N1144), 
        .S1(N1143), .Q(n51979) );
  IMUX40 U57959 ( .A(n51985), .B(n51986), .C(n51987), .D(n51988), .S0(N1144), 
        .S1(N1143), .Q(n51984) );
  MUX41 U57962 ( .A(n51994), .B(n51984), .C(n51989), .D(n51979), .S0(N1146), 
        .S1(N1145), .Q(N6499) );
  IMUX40 U55942 ( .A(n50060), .B(n50061), .C(n50062), .D(n50063), .S0(N1126), 
        .S1(N1125), .Q(n50059) );
  IMUX40 U55943 ( .A(n50065), .B(n50066), .C(n50067), .D(n50068), .S0(N1126), 
        .S1(N1125), .Q(n50064) );
  MUX41 U55946 ( .A(n50074), .B(n50064), .C(n50069), .D(n50059), .S0(N1128), 
        .S1(N1127), .Q(N6362) );
  IMUX40 U49897 ( .A(n44315), .B(n44316), .C(n44317), .D(n44318), .S0(N1072), 
        .S1(n65918), .Q(n44314) );
  IMUX40 U49894 ( .A(n44300), .B(n44301), .C(n44302), .D(n44303), .S0(N1072), 
        .S1(n65917), .Q(n44299) );
  IMUX40 U49895 ( .A(n44305), .B(n44306), .C(n44307), .D(n44308), .S0(N1072), 
        .S1(n65918), .Q(n44304) );
  MUX41 U49898 ( .A(n44314), .B(n44304), .C(n44309), .D(n44299), .S0(N1074), 
        .S1(N1073), .Q(N5964) );
  IMUX40 U61993 ( .A(n55835), .B(n55836), .C(n55837), .D(n55838), .S0(N1180), 
        .S1(n65916), .Q(n55834) );
  IMUX40 U61990 ( .A(n55820), .B(n55821), .C(n55822), .D(n55823), .S0(N1180), 
        .S1(n65918), .Q(n55819) );
  IMUX40 U61991 ( .A(n55825), .B(n55826), .C(n55827), .D(n55828), .S0(N1180), 
        .S1(n65916), .Q(n55824) );
  MUX41 U61994 ( .A(n55834), .B(n55824), .C(n55829), .D(n55819), .S0(N1182), 
        .S1(N1181), .Q(N6777) );
  IMUX40 U64009 ( .A(n57755), .B(n57756), .C(n57757), .D(n57758), .S0(N1198), 
        .S1(N1197), .Q(n57754) );
  IMUX40 U64006 ( .A(n57740), .B(n57741), .C(n57742), .D(n57743), .S0(N1198), 
        .S1(N1197), .Q(n57739) );
  IMUX40 U64007 ( .A(n57745), .B(n57746), .C(n57747), .D(n57748), .S0(N1198), 
        .S1(N1197), .Q(n57744) );
  MUX41 U64010 ( .A(n57754), .B(n57744), .C(n57749), .D(n57739), .S0(N1200), 
        .S1(N1199), .Q(N6914) );
  IMUX40 U16297 ( .A(n12315), .B(n12316), .C(n12317), .D(n12318), .S0(N1060), 
        .S1(N1059), .Q(n12314) );
  IMUX40 U16294 ( .A(n12300), .B(n12301), .C(n12302), .D(n12303), .S0(N1060), 
        .S1(N1059), .Q(n12299) );
  IMUX40 U16295 ( .A(n12305), .B(n12306), .C(n12307), .D(n12308), .S0(N1060), 
        .S1(N1059), .Q(n12304) );
  MUX41 U16298 ( .A(n12314), .B(n12304), .C(n12309), .D(n12299), .S0(N1062), 
        .S1(N1061), .Q(N3599) );
  IMUX40 U18985 ( .A(n14875), .B(n14876), .C(n14877), .D(n14878), .S0(N1084), 
        .S1(N1083), .Q(n14874) );
  IMUX40 U18982 ( .A(n14860), .B(n14861), .C(n14862), .D(n14863), .S0(N1084), 
        .S1(N1083), .Q(n14859) );
  IMUX40 U18983 ( .A(n14865), .B(n14866), .C(n14867), .D(n14868), .S0(N1084), 
        .S1(N1083), .Q(n14864) );
  MUX41 U18986 ( .A(n14874), .B(n14864), .C(n14869), .D(n14859), .S0(N1086), 
        .S1(N1085), .Q(N3758) );
  IMUX40 U31081 ( .A(n26395), .B(n26396), .C(n26397), .D(n26398), .S0(N1192), 
        .S1(N1191), .Q(n26394) );
  IMUX40 U31078 ( .A(n26380), .B(n26381), .C(n26382), .D(n26383), .S0(N1192), 
        .S1(N1191), .Q(n26379) );
  IMUX40 U31079 ( .A(n26385), .B(n26386), .C(n26387), .D(n26388), .S0(N1192), 
        .S1(N1191), .Q(n26384) );
  MUX41 U31082 ( .A(n26394), .B(n26384), .C(n26389), .D(n26379), .S0(N1194), 
        .S1(N1193), .Q(N4571) );
  IMUX40 U33097 ( .A(n28315), .B(n28316), .C(n28317), .D(n28318), .S0(N1210), 
        .S1(n65920), .Q(n28314) );
  IMUX40 U33094 ( .A(n28300), .B(n28301), .C(n28302), .D(n28303), .S0(N1210), 
        .S1(n65919), .Q(n28299) );
  IMUX40 U33095 ( .A(n28305), .B(n28306), .C(n28307), .D(n28308), .S0(N1210), 
        .S1(n65920), .Q(n28304) );
  MUX41 U33098 ( .A(n28314), .B(n28304), .C(n28309), .D(n28299), .S0(N1212), 
        .S1(N1211), .Q(N4708) );
  IMUX40 U53929 ( .A(n48155), .B(n48156), .C(n48157), .D(n48158), .S0(N1108), 
        .S1(N1107), .Q(n48154) );
  IMUX40 U53926 ( .A(n48140), .B(n48141), .C(n48142), .D(n48143), .S0(N1108), 
        .S1(N1107), .Q(n48139) );
  IMUX40 U53927 ( .A(n48145), .B(n48146), .C(n48147), .D(n48148), .S0(N1108), 
        .S1(N1107), .Q(n48144) );
  MUX41 U53930 ( .A(n48154), .B(n48144), .C(n48149), .D(n48139), .S0(N1110), 
        .S1(N1109), .Q(N6226) );
  IMUX40 U14281 ( .A(n10395), .B(n10396), .C(n10397), .D(n10398), .S0(N1042), 
        .S1(N1041), .Q(n10394) );
  IMUX40 U14278 ( .A(n10380), .B(n10381), .C(n10382), .D(n10383), .S0(N1042), 
        .S1(N1041), .Q(n10379) );
  IMUX40 U14279 ( .A(n10385), .B(n10386), .C(n10387), .D(n10388), .S0(N1042), 
        .S1(N1041), .Q(n10384) );
  MUX41 U14282 ( .A(n10394), .B(n10384), .C(n10389), .D(n10379), .S0(N1044), 
        .S1(N1043), .Q(N3472) );
  IMUX40 U35785 ( .A(n30875), .B(n30876), .C(n30877), .D(n30878), .S0(N1234), 
        .S1(N1233), .Q(n30874) );
  IMUX40 U35782 ( .A(n30860), .B(n30861), .C(n30862), .D(n30863), .S0(N1234), 
        .S1(N1233), .Q(n30859) );
  IMUX40 U35783 ( .A(n30865), .B(n30866), .C(n30867), .D(n30868), .S0(N1234), 
        .S1(N1233), .Q(n30864) );
  MUX41 U35786 ( .A(n30874), .B(n30864), .C(n30869), .D(n30859), .S0(N1236), 
        .S1(N1235), .Q(N4920) );
  IMUX40 U41833 ( .A(n36635), .B(n36636), .C(n36637), .D(n36638), .S0(N1000), 
        .S1(N999), .Q(n36634) );
  IMUX40 U41830 ( .A(n36620), .B(n36621), .C(n36622), .D(n36623), .S0(N1000), 
        .S1(N999), .Q(n36619) );
  IMUX40 U41831 ( .A(n36625), .B(n36626), .C(n36627), .D(n36628), .S0(N1000), 
        .S1(N999), .Q(n36624) );
  MUX41 U41834 ( .A(n36634), .B(n36624), .C(n36629), .D(n36619), .S0(N1002), 
        .S1(N1001), .Q(N5400) );
  IMUX40 U43849 ( .A(n38555), .B(n38556), .C(n38557), .D(n38558), .S0(N1018), 
        .S1(N1017), .Q(n38554) );
  IMUX40 U43846 ( .A(n38540), .B(n38541), .C(n38542), .D(n38543), .S0(N1018), 
        .S1(N1017), .Q(n38539) );
  IMUX40 U43847 ( .A(n38545), .B(n38546), .C(n38547), .D(n38548), .S0(N1018), 
        .S1(N1017), .Q(n38544) );
  MUX41 U43850 ( .A(n38554), .B(n38544), .C(n38549), .D(n38539), .S0(N1020), 
        .S1(N1019), .Q(N5555) );
  IMUX40 U45865 ( .A(n40475), .B(n40476), .C(n40477), .D(n40478), .S0(N1036), 
        .S1(N1035), .Q(n40474) );
  IMUX40 U45862 ( .A(n40460), .B(n40461), .C(n40462), .D(n40463), .S0(N1036), 
        .S1(N1035), .Q(n40459) );
  IMUX40 U45863 ( .A(n40465), .B(n40466), .C(n40467), .D(n40468), .S0(N1036), 
        .S1(N1035), .Q(n40464) );
  MUX41 U45866 ( .A(n40474), .B(n40464), .C(n40469), .D(n40459), .S0(N1038), 
        .S1(N1037), .Q(N5710) );
  IMUX40 U68041 ( .A(n61595), .B(n61596), .C(n61597), .D(n61598), .S0(N1234), 
        .S1(N1233), .Q(n61594) );
  IMUX40 U68038 ( .A(n61580), .B(n61581), .C(n61582), .D(n61583), .S0(N1234), 
        .S1(N1233), .Q(n61579) );
  IMUX40 U68039 ( .A(n61585), .B(n61586), .C(n61587), .D(n61588), .S0(N1234), 
        .S1(N1233), .Q(n61584) );
  MUX41 U68042 ( .A(n61594), .B(n61584), .C(n61589), .D(n61579), .S0(N1236), 
        .S1(N1235), .Q(N7190) );
  IMUX40 U22345 ( .A(n18075), .B(n18076), .C(n18077), .D(n18078), .S0(N1114), 
        .S1(N1113), .Q(n18074) );
  IMUX40 U22342 ( .A(n18060), .B(n18061), .C(n18062), .D(n18063), .S0(N1114), 
        .S1(N1113), .Q(n18059) );
  IMUX40 U22343 ( .A(n18065), .B(n18066), .C(n18067), .D(n18068), .S0(N1114), 
        .S1(N1113), .Q(n18064) );
  MUX41 U22346 ( .A(n18074), .B(n18064), .C(n18069), .D(n18059), .S0(N1116), 
        .S1(N1115), .Q(N3988) );
  IMUX40 U23689 ( .A(n19355), .B(n19356), .C(n19357), .D(n19358), .S0(N838), 
        .S1(N837), .Q(n19354) );
  IMUX40 U23686 ( .A(n19340), .B(n19341), .C(n19342), .D(n19343), .S0(N838), 
        .S1(N837), .Q(n19339) );
  IMUX40 U23687 ( .A(n19345), .B(n19346), .C(n19347), .D(n19348), .S0(N838), 
        .S1(N837), .Q(n19344) );
  MUX41 U23690 ( .A(n19354), .B(n19344), .C(n19349), .D(n19339), .S0(N840), 
        .S1(N839), .Q(N4092) );
  IMUX40 U38473 ( .A(n33435), .B(n33436), .C(n33437), .D(n33438), .S0(N970), 
        .S1(N969), .Q(n33434) );
  IMUX40 U38470 ( .A(n33420), .B(n33421), .C(n33422), .D(n33423), .S0(N970), 
        .S1(N969), .Q(n33419) );
  IMUX40 U38471 ( .A(n33425), .B(n33426), .C(n33427), .D(n33428), .S0(N970), 
        .S1(N969), .Q(n33424) );
  MUX41 U38474 ( .A(n33434), .B(n33424), .C(n33429), .D(n33419), .S0(N972), 
        .S1(N971), .Q(N5090) );
  IMUX40 U24361 ( .A(n19995), .B(n19996), .C(n19997), .D(n19998), .S0(N844), 
        .S1(N843), .Q(n19994) );
  IMUX40 U24358 ( .A(n19980), .B(n19981), .C(n19982), .D(n19983), .S0(N844), 
        .S1(N843), .Q(n19979) );
  IMUX40 U24359 ( .A(n19985), .B(n19986), .C(n19987), .D(n19988), .S0(N844), 
        .S1(N843), .Q(n19984) );
  MUX41 U24362 ( .A(n19994), .B(n19984), .C(n19989), .D(n19979), .S0(N846), 
        .S1(N845), .Q(N4124) );
  IMUX40 U10246 ( .A(n6540), .B(n6541), .C(n6542), .D(n6543), .S0(N718), .S1(
        N717), .Q(n6539) );
  IMUX40 U10247 ( .A(n6545), .B(n6546), .C(n6547), .D(n6548), .S0(N718), .S1(
        N717), .Q(n6544) );
  IMUX40 U18313 ( .A(n14235), .B(n14236), .C(n14237), .D(n14238), .S0(N1078), 
        .S1(N1077), .Q(n14234) );
  IMUX40 U18310 ( .A(n14220), .B(n14221), .C(n14222), .D(n14223), .S0(N1078), 
        .S1(N1077), .Q(n14219) );
  IMUX40 U18311 ( .A(n14225), .B(n14226), .C(n14227), .D(n14228), .S0(N1078), 
        .S1(N1077), .Q(n14224) );
  IMUX40 U17641 ( .A(n13595), .B(n13596), .C(n13597), .D(n13598), .S0(N1072), 
        .S1(n65918), .Q(n13594) );
  IMUX40 U17638 ( .A(n13580), .B(n13581), .C(n13582), .D(n13583), .S0(N1072), 
        .S1(n65918), .Q(n13579) );
  IMUX40 U17639 ( .A(n13585), .B(n13586), .C(n13587), .D(n13588), .S0(N1072), 
        .S1(n65918), .Q(n13584) );
  IMUX40 U29737 ( .A(n25115), .B(n25116), .C(n25117), .D(n25118), .S0(N1180), 
        .S1(n65916), .Q(n25114) );
  IMUX40 U29734 ( .A(n25100), .B(n25101), .C(n25102), .D(n25103), .S0(N1180), 
        .S1(n65916), .Q(n25099) );
  IMUX40 U29735 ( .A(n25105), .B(n25106), .C(n25107), .D(n25108), .S0(N1180), 
        .S1(n65915), .Q(n25104) );
  IMUX40 U32425 ( .A(n27675), .B(n27676), .C(n27677), .D(n27678), .S0(N1204), 
        .S1(N1203), .Q(n27674) );
  IMUX40 U32422 ( .A(n27660), .B(n27661), .C(n27662), .D(n27663), .S0(N1204), 
        .S1(N1203), .Q(n27659) );
  IMUX40 U32423 ( .A(n27665), .B(n27666), .C(n27667), .D(n27668), .S0(N1204), 
        .S1(N1203), .Q(n27664) );
  IMUX40 U31753 ( .A(n27035), .B(n27036), .C(n27037), .D(n27038), .S0(N1198), 
        .S1(N1197), .Q(n27034) );
  IMUX40 U31750 ( .A(n27020), .B(n27021), .C(n27022), .D(n27023), .S0(N1198), 
        .S1(N1197), .Q(n27019) );
  IMUX40 U31751 ( .A(n27025), .B(n27026), .C(n27027), .D(n27028), .S0(N1198), 
        .S1(N1197), .Q(n27024) );
  IMUX40 U9577 ( .A(n5915), .B(n5916), .C(n5917), .D(n5918), .S0(N1000), .S1(
        N999), .Q(n5914) );
  IMUX40 U9574 ( .A(n5900), .B(n5901), .C(n5902), .D(n5903), .S0(N1000), .S1(
        N999), .Q(n5899) );
  IMUX40 U9575 ( .A(n5905), .B(n5906), .C(n5907), .D(n5908), .S0(N1000), .S1(
        N999), .Q(n5904) );
  IMUX40 U12265 ( .A(n8475), .B(n8476), .C(n8477), .D(n8478), .S0(N1024), .S1(
        N1023), .Q(n8474) );
  IMUX40 U12262 ( .A(n8460), .B(n8461), .C(n8462), .D(n8463), .S0(N1024), .S1(
        N1023), .Q(n8459) );
  IMUX40 U12263 ( .A(n8465), .B(n8466), .C(n8467), .D(n8468), .S0(N1024), .S1(
        N1023), .Q(n8464) );
  MUX41 U12266 ( .A(n8474), .B(n8464), .C(n8469), .D(n8459), .S0(N1026), .S1(
        N1025), .Q(N3317) );
  IMUX40 U11593 ( .A(n7835), .B(n7836), .C(n7837), .D(n7838), .S0(N1018), .S1(
        N1017), .Q(n7834) );
  IMUX40 U11590 ( .A(n7820), .B(n7821), .C(n7822), .D(n7823), .S0(N1018), .S1(
        N1017), .Q(n7819) );
  IMUX40 U11591 ( .A(n7825), .B(n7826), .C(n7827), .D(n7828), .S0(N1018), .S1(
        N1017), .Q(n7824) );
  MUX41 U11594 ( .A(n7834), .B(n7824), .C(n7829), .D(n7819), .S0(N1020), .S1(
        N1019), .Q(N3285) );
  IMUX40 U13609 ( .A(n9755), .B(n9756), .C(n9757), .D(n9758), .S0(N1036), .S1(
        N1035), .Q(n9754) );
  IMUX40 U13606 ( .A(n9740), .B(n9741), .C(n9742), .D(n9743), .S0(N1036), .S1(
        N1035), .Q(n9739) );
  IMUX40 U13607 ( .A(n9745), .B(n9746), .C(n9747), .D(n9748), .S0(N1036), .S1(
        N1035), .Q(n9744) );
  IMUX40 U30409 ( .A(n25755), .B(n25756), .C(n25757), .D(n25758), .S0(N1186), 
        .S1(N1185), .Q(n25754) );
  IMUX40 U30406 ( .A(n25740), .B(n25741), .C(n25742), .D(n25743), .S0(N1186), 
        .S1(N1185), .Q(n25739) );
  IMUX40 U30407 ( .A(n25745), .B(n25746), .C(n25747), .D(n25748), .S0(N1186), 
        .S1(N1185), .Q(n25744) );
  IMUX40 U55273 ( .A(n49435), .B(n49436), .C(n49437), .D(n49438), .S0(N1120), 
        .S1(n65917), .Q(n49434) );
  IMUX40 U55270 ( .A(n49420), .B(n49421), .C(n49422), .D(n49423), .S0(N1120), 
        .S1(n65917), .Q(n49419) );
  IMUX40 U55271 ( .A(n49425), .B(n49426), .C(n49427), .D(n49428), .S0(N11412), 
        .S1(n65917), .Q(n49424) );
  MUX41 U55274 ( .A(n49434), .B(n49424), .C(n49429), .D(n49419), .S0(N1122), 
        .S1(N1121), .Q(N6290) );
  IMUX40 U37128 ( .A(n32150), .B(n32151), .C(n32152), .D(n32153), .S0(N958), 
        .S1(N957), .Q(n32149) );
  IMUX40 U37126 ( .A(n32140), .B(n32141), .C(n32142), .D(n32143), .S0(N958), 
        .S1(N957), .Q(n32139) );
  IMUX40 U37127 ( .A(n32145), .B(n32146), .C(n32147), .D(n32148), .S0(N958), 
        .S1(N957), .Q(n32144) );
  MUX41 U37130 ( .A(n32154), .B(n32144), .C(n32149), .D(n32139), .S0(N960), 
        .S1(N959), .Q(N4984) );
  IMUX40 U69384 ( .A(n62870), .B(n62871), .C(n62872), .D(n62873), .S0(N1246), 
        .S1(N1245), .Q(n62869) );
  IMUX40 U69382 ( .A(n62860), .B(n62861), .C(n62862), .D(n62863), .S0(N1246), 
        .S1(N1245), .Q(n62859) );
  IMUX40 U69383 ( .A(n62865), .B(n62866), .C(n62867), .D(n62868), .S0(N1246), 
        .S1(N1245), .Q(n62864) );
  MUX41 U69386 ( .A(n62874), .B(n62864), .C(n62869), .D(n62859), .S0(N1248), 
        .S1(N1247), .Q(N7254) );
  IMUX40 U41158 ( .A(n35980), .B(n35981), .C(n35982), .D(n35983), .S0(N994), 
        .S1(N993), .Q(n35979) );
  IMUX40 U41159 ( .A(n35985), .B(n35986), .C(n35987), .D(n35988), .S0(N994), 
        .S1(N993), .Q(n35984) );
  MUX41 U41162 ( .A(n35994), .B(n35984), .C(n35989), .D(n35979), .S0(N996), 
        .S1(N995), .Q(N5310) );
  IMUX40 U43174 ( .A(n37900), .B(n37901), .C(n37902), .D(n37903), .S0(N1012), 
        .S1(N1011), .Q(n37899) );
  IMUX40 U43175 ( .A(n37905), .B(n37906), .C(n37907), .D(n37908), .S0(N1012), 
        .S1(N1011), .Q(n37904) );
  MUX41 U43178 ( .A(n37914), .B(n37904), .C(n37909), .D(n37899), .S0(N1014), 
        .S1(N1013), .Q(N5464) );
  IMUX40 U45190 ( .A(n39820), .B(n39821), .C(n39822), .D(n39823), .S0(N1030), 
        .S1(N1029), .Q(n39819) );
  IMUX40 U45191 ( .A(n39825), .B(n39826), .C(n39827), .D(n39828), .S0(N1030), 
        .S1(N1029), .Q(n39824) );
  MUX41 U45194 ( .A(n39834), .B(n39824), .C(n39829), .D(n39819), .S0(N1032), 
        .S1(N1031), .Q(N5619) );
  IMUX40 U71398 ( .A(n64780), .B(n64781), .C(n64782), .D(n64783), .S0(N1264), 
        .S1(N1263), .Q(n64779) );
  IMUX40 U71399 ( .A(n64785), .B(n64786), .C(n64787), .D(n64788), .S0(N1264), 
        .S1(N1263), .Q(n64784) );
  MUX41 U71402 ( .A(n64794), .B(n64784), .C(n64789), .D(n64779), .S0(N1266), 
        .S1(N1265), .Q(N7392) );
  IMUX40 U57286 ( .A(n51340), .B(n51341), .C(n51342), .D(n51343), .S0(N1138), 
        .S1(n65919), .Q(n51339) );
  IMUX40 U57287 ( .A(n51345), .B(n51346), .C(n51347), .D(n51348), .S0(N1138), 
        .S1(n65919), .Q(n51344) );
  MUX41 U57290 ( .A(n51354), .B(n51344), .C(n51349), .D(n51339), .S0(N1140), 
        .S1(N1139), .Q(N6426) );
  IMUX40 U49225 ( .A(n43675), .B(n43676), .C(n43677), .D(n43678), .S0(N1066), 
        .S1(n65920), .Q(n43674) );
  IMUX40 U49222 ( .A(n43660), .B(n43661), .C(n43662), .D(n43663), .S0(N1066), 
        .S1(n65920), .Q(n43659) );
  IMUX40 U49223 ( .A(n43665), .B(n43666), .C(n43667), .D(n43668), .S0(N1066), 
        .S1(n65920), .Q(n43664) );
  MUX41 U49226 ( .A(n43674), .B(n43664), .C(n43669), .D(n43659), .S0(N1068), 
        .S1(N1067), .Q(N5901) );
  IMUX40 U51241 ( .A(n45595), .B(n45596), .C(n45597), .D(n45598), .S0(N1084), 
        .S1(N1083), .Q(n45594) );
  IMUX40 U51238 ( .A(n45580), .B(n45581), .C(n45582), .D(n45583), .S0(N1084), 
        .S1(N1083), .Q(n45579) );
  IMUX40 U51239 ( .A(n45585), .B(n45586), .C(n45587), .D(n45588), .S0(N1084), 
        .S1(N1083), .Q(n45584) );
  MUX41 U51242 ( .A(n45594), .B(n45584), .C(n45589), .D(n45579), .S0(N1086), 
        .S1(N1085), .Q(N6028) );
  IMUX40 U63337 ( .A(n57115), .B(n57116), .C(n57117), .D(n57118), .S0(N1192), 
        .S1(N1191), .Q(n57114) );
  IMUX40 U63334 ( .A(n57100), .B(n57101), .C(n57102), .D(n57103), .S0(N1192), 
        .S1(N1191), .Q(n57099) );
  IMUX40 U63335 ( .A(n57105), .B(n57106), .C(n57107), .D(n57108), .S0(N1192), 
        .S1(N1191), .Q(n57104) );
  MUX41 U63338 ( .A(n57114), .B(n57104), .C(n57109), .D(n57099), .S0(N1194), 
        .S1(N1193), .Q(N6841) );
  IMUX40 U65353 ( .A(n59035), .B(n59036), .C(n59037), .D(n59038), .S0(N1210), 
        .S1(n65920), .Q(n59034) );
  IMUX40 U65350 ( .A(n59020), .B(n59021), .C(n59022), .D(n59023), .S0(N1210), 
        .S1(n65919), .Q(n59019) );
  IMUX40 U65351 ( .A(n59025), .B(n59026), .C(n59027), .D(n59028), .S0(N1210), 
        .S1(n65919), .Q(n59024) );
  MUX41 U65354 ( .A(n59034), .B(n59024), .C(n59029), .D(n59019), .S0(N1212), 
        .S1(N1211), .Q(N6978) );
  IMUX40 U27049 ( .A(n22555), .B(n22556), .C(n22557), .D(n22558), .S0(N1156), 
        .S1(n65917), .Q(n22554) );
  IMUX40 U27046 ( .A(n22540), .B(n22541), .C(n22542), .D(n22543), .S0(N1156), 
        .S1(n65918), .Q(n22539) );
  IMUX40 U27047 ( .A(n22545), .B(n22546), .C(n22547), .D(n22548), .S0(N1156), 
        .S1(n65918), .Q(n22544) );
  MUX41 U27050 ( .A(n22554), .B(n22544), .C(n22549), .D(n22539), .S0(N1158), 
        .S1(N1157), .Q(N4293) );
  IMUX40 U47209 ( .A(n41755), .B(n41756), .C(n41757), .D(n41758), .S0(N1048), 
        .S1(N1047), .Q(n41754) );
  IMUX40 U47206 ( .A(n41740), .B(n41741), .C(n41742), .D(n41743), .S0(N1048), 
        .S1(N1047), .Q(n41739) );
  IMUX40 U47207 ( .A(n41745), .B(n41746), .C(n41747), .D(n41748), .S0(N1048), 
        .S1(N1047), .Q(n41744) );
  MUX41 U47210 ( .A(n41754), .B(n41744), .C(n41749), .D(n41739), .S0(N1050), 
        .S1(N1049), .Q(N5774) );
  IMUX40 U59305 ( .A(n53275), .B(n53276), .C(n53277), .D(n53278), .S0(N1156), 
        .S1(n65918), .Q(n53274) );
  IMUX40 U59302 ( .A(n53260), .B(n53261), .C(n53262), .D(n53263), .S0(N1156), 
        .S1(n65917), .Q(n53259) );
  IMUX40 U59303 ( .A(n53265), .B(n53266), .C(n53267), .D(n53268), .S0(N1156), 
        .S1(n65918), .Q(n53264) );
  MUX41 U59306 ( .A(n53274), .B(n53264), .C(n53269), .D(n53259), .S0(N1158), 
        .S1(N1157), .Q(N6563) );
  IMUX40 U29065 ( .A(n24475), .B(n24476), .C(n24477), .D(n24478), .S0(N1174), 
        .S1(N1173), .Q(n24474) );
  IMUX40 U29062 ( .A(n24460), .B(n24461), .C(n24462), .D(n24463), .S0(N1174), 
        .S1(N1173), .Q(n24459) );
  IMUX40 U29063 ( .A(n24465), .B(n24466), .C(n24467), .D(n24468), .S0(N1174), 
        .S1(N1173), .Q(n24464) );
  MUX41 U29066 ( .A(n24474), .B(n24464), .C(n24469), .D(n24459), .S0(N1176), 
        .S1(N1175), .Q(N4432) );
  IMUX40 U61321 ( .A(n55195), .B(n55196), .C(n55197), .D(n55198), .S0(N1174), 
        .S1(N1173), .Q(n55194) );
  IMUX40 U61318 ( .A(n55180), .B(n55181), .C(n55182), .D(n55183), .S0(N1174), 
        .S1(N1173), .Q(n55179) );
  IMUX40 U61319 ( .A(n55185), .B(n55186), .C(n55187), .D(n55188), .S0(N1174), 
        .S1(N1173), .Q(n55184) );
  MUX41 U61322 ( .A(n55194), .B(n55184), .C(n55189), .D(n55179), .S0(N1176), 
        .S1(N1175), .Q(N6702) );
  MUX41 U54602 ( .A(n48794), .B(n48784), .C(n48789), .D(n48779), .S0(N1116), 
        .S1(N1115), .Q(N6258) );
  MUX41 U33770 ( .A(n28954), .B(n28944), .C(n28949), .D(n28939), .S0(N1218), 
        .S1(N1217), .Q(N4781) );
  MUX41 U34442 ( .A(n29594), .B(n29584), .C(n29589), .D(n29579), .S0(N1224), 
        .S1(N1223), .Q(N4813) );
  MUX41 U66026 ( .A(n59674), .B(n59664), .C(n59669), .D(n59659), .S0(N1218), 
        .S1(N1217), .Q(N7051) );
  MUX41 U66698 ( .A(n60314), .B(n60304), .C(n60309), .D(n60299), .S0(N1224), 
        .S1(N1223), .Q(N7083) );
  MUX41 U47882 ( .A(n42394), .B(n42384), .C(n42389), .D(n42379), .S0(N1056), 
        .S1(N1055), .Q(N5837) );
  MUX41 U48554 ( .A(n43034), .B(n43024), .C(n43029), .D(n43019), .S0(N1062), 
        .S1(N1061), .Q(N5869) );
  MUX41 U50570 ( .A(n44954), .B(n44944), .C(n44949), .D(n44939), .S0(N1080), 
        .S1(N1079), .Q(N5996) );
  DF1 \O_play_reg[3]  ( .D(O[3]), .C(CLK), .Q(O_play[3]) );
  DF1 \O_play_reg[2]  ( .D(O[2]), .C(CLK), .Q(O_play[2]) );
  DF1 \O_play_reg[1]  ( .D(O[1]), .C(CLK), .Q(O_play[1]) );
  DF1 \G_play_reg[2]  ( .D(G[2]), .C(CLK), .Q(G_play[2]) );
  DF1 \G_play_reg[1]  ( .D(G[1]), .C(CLK), .Q(G_play[1]) );
  IMUX21 U7175 ( .A(n3725), .B(n3726), .S(n65946), .Q(N1362) );
  IMUX21 U7176 ( .A(n3727), .B(n3728), .S(n65946), .Q(N1361) );
  IMUX21 U7178 ( .A(n3731), .B(n3732), .S(n65946), .Q(N1359) );
  IMUX21 U7370 ( .A(n3859), .B(n3860), .S(n65936), .Q(N1902) );
  IMUX21 U7177 ( .A(n3729), .B(n3730), .S(n65946), .Q(N1360) );
  IMUX21 U7369 ( .A(n3857), .B(n3858), .S(n65936), .Q(N1903) );
  DF3 \O_play_reg[0]  ( .D(O[0]), .C(CLK), .Q(n65419), .QN(n65740) );
  DF3 \G_play_reg[0]  ( .D(G[0]), .C(CLK), .Q(n65420), .QN(n65742) );
  CLKIN6 U72070 ( .A(m[3]), .Q(n66739) );
  CLKIN6 U72071 ( .A(m[3]), .Q(n66684) );
  CLKIN6 U72072 ( .A(m[3]), .Q(N3196) );
  NOR31 U72073 ( .A(n65609), .B(n65544), .C(m[3]), .Q(n66728) );
  OAI222 U72074 ( .A(n65610), .B(m[3]), .C(n65604), .D(m[3]), .Q(N4709) );
  OAI222 U72075 ( .A(n65610), .B(m[3]), .C(n65604), .D(m[3]), .Q(N3505) );
  CLKIN6 U72076 ( .A(m[3]), .Q(N4986) );
  CLKIN6 U72077 ( .A(m[3]), .Q(n66824) );
  NOR31 U72078 ( .A(n65609), .B(n65544), .C(m[3]), .Q(n66683) );
  NOR31 U72079 ( .A(n65609), .B(n65544), .C(m[3]), .Q(n66846) );
  OAI222 U72080 ( .A(n65610), .B(m[3]), .C(n65604), .D(m[3]), .Q(N4572) );
  CLKIN6 U72081 ( .A(m[3]), .Q(N4295) );
  CLKIN6 U72082 ( .A(m[3]), .Q(n66687) );
  NOR40 U72083 ( .A(n65544), .B(m[3]), .C(n65610), .D(n65604), .Q(n66686) );
  INV3 U72084 ( .A(n65990), .Q(\add_1_root_add_0_root_sub_328_4_cf/carry[4] )
         );
  INV3 U72085 ( .A(n66057), .Q(\r12188/carry [4]) );
  INV3 U72086 ( .A(n65988), .Q(\add_1_root_add_0_root_sub_331_4_cf/carry[4] )
         );
  INV3 U72087 ( .A(n66035), .Q(\add_1_root_add_0_root_sub_397_8_cf/carry[4] )
         );
  XOR21 U72088 ( .A(n65758), .B(n65905), .Q(N1130) );
  XOR21 U72089 ( .A(n65758), .B(n65909), .Q(N1148) );
  ADD22 U72090 ( .A(n65758), .B(n65841), .CO(\r31196/carry [2]), .S(N1172) );
  ADD22 U72091 ( .A(n65758), .B(n65842), .CO(\r32997/carry [2]), .S(N1184) );
  XOR21 U72092 ( .A(n65594), .B(n65585), .Q(N11412) );
  INV3 U72093 ( .A(n65985), .Q(\add_1_root_add_0_root_sub_348_9_cf/carry [4])
         );
  XNR21 U72094 ( .A(n65605), .B(n65583), .Q(N4602) );
  AOI211 U72095 ( .A(n3676), .B(n66567), .C(n3274), .Q(n3325) );
  AOI211 U72096 ( .A(n66567), .B(n3655), .C(n3274), .Q(n3355) );
  OAI212 U72097 ( .A(n65817), .B(n65770), .C(n66103), .Q(N1046) );
  OAI212 U72098 ( .A(n65817), .B(n65775), .C(n66097), .Q(N1034) );
  OAI212 U72099 ( .A(n65809), .B(n65773), .C(n66114), .Q(N1040) );
  INV3 U72100 ( .A(n66018), .Q(\r34786/carry [3]) );
  INV3 U72101 ( .A(n66027), .Q(\r38360/carry [4]) );
  INV3 U72102 ( .A(n66008), .Q(\r32996/carry [4]) );
  INV3 U72103 ( .A(n65993), .Q(\add_1_root_add_0_root_sub_328_8_cf/carry[2] )
         );
  INV3 U72104 ( .A(n65986), .Q(\add_1_root_add_0_root_sub_348_9_cf/carry [3])
         );
  INV3 U72105 ( .A(n66010), .Q(\r41369/carry[4] ) );
  IMUX40 U72106 ( .A(n14234), .B(n14224), .C(n14229), .D(n14219), .S0(N1080), 
        .S1(N1079), .Q(n65421) );
  IMUX40 U72107 ( .A(n27674), .B(n27664), .C(n27669), .D(n27659), .S0(N1206), 
        .S1(N1205), .Q(n65422) );
  IMUX40 U72108 ( .A(n25754), .B(n25744), .C(n25749), .D(n25739), .S0(N1188), 
        .S1(N1187), .Q(n65423) );
  IMUX40 U72109 ( .A(n6554), .B(n6544), .C(n6549), .D(n6539), .S0(N720), .S1(
        N719), .Q(n65424) );
  NAND22 U72110 ( .A(n66082), .B(n66083), .Q(N1946) );
  NAND22 U72111 ( .A(n66108), .B(\sub_140_b0/carry [5]), .Q(n65963) );
  NAND22 U72112 ( .A(n66122), .B(\sub_171_b0/carry [5]), .Q(n65976) );
  AOI211 U72113 ( .A(n65740), .B(N1836), .C(n66872), .Q(n66871) );
  IMUX40 U72114 ( .A(n13594), .B(n13584), .C(n13589), .D(n13579), .S0(N1074), 
        .S1(N1073), .Q(n65425) );
  IMUX40 U72115 ( .A(n27034), .B(n27024), .C(n27029), .D(n27019), .S0(N1200), 
        .S1(N1199), .Q(n65426) );
  IMUX40 U72116 ( .A(n25114), .B(n25104), .C(n25109), .D(n25099), .S0(N1182), 
        .S1(N1181), .Q(n65427) );
  IMUX40 U72117 ( .A(n5914), .B(n5904), .C(n5909), .D(n5899), .S0(N1002), .S1(
        N1001), .Q(n65428) );
  IMUX40 U72118 ( .A(n11674), .B(n11664), .C(n11669), .D(n11659), .S0(N1056), 
        .S1(N1055), .Q(n65429) );
  IMUX40 U72119 ( .A(n17434), .B(n17424), .C(n17429), .D(n17419), .S0(N1110), 
        .S1(N1109), .Q(n65430) );
  IMUX40 U72120 ( .A(n3994), .B(n3984), .C(n3989), .D(n3979), .S0(N696), .S1(
        N695), .Q(n65431) );
  IMUX40 U72121 ( .A(n9754), .B(n9744), .C(n9749), .D(n9739), .S0(N1038), .S1(
        N1037), .Q(n65432) );
  CLKIN0 U72122 ( .A(n3721), .Q(n65433) );
  INV3 U72123 ( .A(n65433), .Q(n65434) );
  OAI210 U72124 ( .A(n1683), .B(n1681), .C(n1684), .Q(n3721) );
  CLKIN0 U72125 ( .A(n3722), .Q(n65435) );
  INV3 U72126 ( .A(n65435), .Q(n65436) );
  OAI210 U72127 ( .A(n1683), .B(n1682), .C(n1723), .Q(n3722) );
  XOR22 U72128 ( .A(N3382), .B(n65584), .Q(N1042) );
  XOR22 U72129 ( .A(N3209), .B(n65582), .Q(N1018) );
  XOR22 U72130 ( .A(N11268), .B(n65585), .Q(N1066) );
  XOR22 U72131 ( .A(N11292), .B(n65581), .Q(N1084) );
  XOR22 U72132 ( .A(N11262), .B(n65583), .Q(N1060) );
  XOR22 U72133 ( .A(n[3]), .B(N3200), .Q(N1180) );
  XOR22 U72134 ( .A(N11286), .B(n65583), .Q(N1078) );
  XOR22 U72135 ( .A(n65594), .B(n65578), .Q(N1156) );
  XOR22 U72136 ( .A(N11466), .B(n65581), .Q(N1204) );
  XOR22 U72137 ( .A(N11496), .B(n65582), .Q(N1222) );
  XOR22 U72138 ( .A(N3054), .B(n65578), .Q(N1000) );
  XOR22 U72139 ( .A(N3364), .B(N3200), .Q(N1036) );
  XOR22 U72140 ( .A(N3400), .B(n65579), .Q(N1048) );
  XOR22 U72141 ( .A(N3227), .B(n65578), .Q(N1024) );
  XOR22 U72142 ( .A(N11460), .B(N3200), .Q(N1198) );
  XOR22 U72143 ( .A(N11472), .B(n65579), .Q(N1210) );
  XOR22 U72144 ( .A(N11514), .B(N3200), .Q(N1234) );
  XOR22 U72145 ( .A(N11256), .B(n65585), .Q(N1054) );
  XOR22 U72146 ( .A(N11490), .B(n65579), .Q(N1216) );
  XOR22 U72147 ( .A(n65594), .B(n65580), .Q(N1072) );
  XOR22 U72148 ( .A(n65594), .B(n65578), .Q(N1168) );
  XOR22 U72149 ( .A(N11436), .B(N3200), .Q(N1192) );
  XOR22 U72150 ( .A(N11322), .B(n65585), .Q(N1108) );
  XOR20 U72151 ( .A(n65918), .B(n65758), .Q(N975) );
  XNR20 U72152 ( .A(n65755), .B(n65891), .Q(N692) );
  XNR20 U72153 ( .A(n65754), .B(n65894), .Q(N698) );
  XOR20 U72154 ( .A(n65758), .B(n65903), .Q(N860) );
  XNR20 U72155 ( .A(n65758), .B(n65866), .Q(n65438) );
  XNR20 U72156 ( .A(n65905), .B(n65758), .Q(n65437) );
  XNR21 U72157 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65918), 
        .Q(N1221) );
  XNR21 U72158 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65918), 
        .Q(N1203) );
  XNR21 U72159 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65918), 
        .Q(N1059) );
  XNR21 U72160 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65918), 
        .Q(N1083) );
  XNR21 U72161 ( .A(n65748), .B(N1167), .Q(N1215) );
  XNR21 U72162 ( .A(n65758), .B(n65918), .Q(N1053) );
  XNR21 U72163 ( .A(n65758), .B(n65918), .Q(N1077) );
  XNR21 U72164 ( .A(n65747), .B(n65917), .Q(N1233) );
  XNR21 U72165 ( .A(n65750), .B(n65916), .Q(N1197) );
  XOR21 U72166 ( .A(n65915), .B(n65758), .Q(N1107) );
  XOR21 U72167 ( .A(N1167), .B(n65758), .Q(N1191) );
  XOR21 U72168 ( .A(N11544), .B(n65579), .Q(N976) );
  XOR21 U72169 ( .A(N11532), .B(N3200), .Q(N1264) );
  XOR21 U72170 ( .A(N11346), .B(n65579), .Q(N1138) );
  XOR21 U72171 ( .A(N11334), .B(n65578), .Q(N1126) );
  XOR21 U72172 ( .A(N11370), .B(N3200), .Q(N1144) );
  XOR21 U72173 ( .A(N11394), .B(n65579), .Q(N1162) );
  XOR21 U72174 ( .A(N11382), .B(N3200), .Q(N856) );
  XOR21 U72175 ( .A(N11406), .B(n65579), .Q(N874) );
  XOR21 U72176 ( .A(n65594), .B(n65577), .Q(N1240) );
  XOR21 U72177 ( .A(N5170), .B(n65578), .Q(N982) );
  XOR21 U72178 ( .A(N3245), .B(N3200), .Q(N742) );
  XOR21 U72179 ( .A(N5515), .B(n65578), .Q(N1030) );
  XOR21 U72180 ( .A(N5342), .B(n65578), .Q(N1006) );
  XOR21 U72181 ( .A(N5206), .B(n65578), .Q(N994) );
  XOR21 U72182 ( .A(N3072), .B(n65579), .Q(N718) );
  XOR21 U72183 ( .A(N2936), .B(n65578), .Q(N706) );
  XOR21 U72184 ( .A(n[3]), .B(n65577), .Q(N952) );
  XOR21 U72185 ( .A(n[3]), .B(N3200), .Q(N964) );
  XOR21 U72186 ( .A(n[3]), .B(n65579), .Q(N1252) );
  XOR21 U72187 ( .A(n[3]), .B(n65578), .Q(N1228) );
  XOR21 U72188 ( .A(n[3]), .B(n65578), .Q(N940) );
  XOR21 U72189 ( .A(n66104), .B(n65532), .Q(N11206) );
  XNR21 U72190 ( .A(n65917), .B(n65758), .Q(N837) );
  XNR21 U72191 ( .A(n65758), .B(n65916), .Q(N1125) );
  XNR21 U72192 ( .A(n65758), .B(N1167), .Q(N1143) );
  XNR21 U72193 ( .A(n65758), .B(n65915), .Q(N1161) );
  XNR21 U72194 ( .A(n65751), .B(n65918), .Q(N855) );
  XNR21 U72195 ( .A(n65749), .B(n65918), .Q(N873) );
  XNR21 U72196 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65917), 
        .Q(N1131) );
  XNR21 U72197 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65915), 
        .Q(N1149) );
  XNR21 U72198 ( .A(N1167), .B(\add_0_root_add_0_root_sub_325_8_cf/carry [2]), 
        .Q(N843) );
  XNR21 U72199 ( .A(n65916), .B(n66114), .Q(N693) );
  XNR21 U72200 ( .A(n65915), .B(n66103), .Q(N699) );
  XNR21 U72201 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65918), 
        .Q(N861) );
  XOR21 U72202 ( .A(N11340), .B(n65584), .Q(N1132) );
  XOR21 U72203 ( .A(N11376), .B(n65582), .Q(N1150) );
  XOR21 U72204 ( .A(N11388), .B(n65584), .Q(N862) );
  XOR21 U72205 ( .A(N5188), .B(n65584), .Q(N988) );
  XOR21 U72206 ( .A(N5360), .B(n65581), .Q(N1012) );
  XOR21 U72207 ( .A(N3090), .B(n65585), .Q(N724) );
  XOR31 U72208 ( .A(n[5]), .B(N11362), .C(
        \add_0_root_add_0_root_sub_325_12_cf/carry [5]), .Q(N852) );
  XOR31 U72209 ( .A(N3900), .B(n[5]), .C(\r13449/carry[5] ), .Q(N1122) );
  XOR31 U72210 ( .A(N3638), .B(n[5]), .C(\r12187/carry[5] ), .Q(N1074) );
  XOR31 U72211 ( .A(N3511), .B(N11260), .C(\r11557/carry [5]), .Q(N1062) );
  XOR31 U72212 ( .A(N3511), .B(N11254), .C(\r11556/carry [5]), .Q(N1056) );
  XOR31 U72213 ( .A(N3638), .B(N11290), .C(\r12191/carry [5]), .Q(N1086) );
  XOR31 U72214 ( .A(N3511), .B(N11266), .C(\r11558/carry [5]), .Q(N1068) );
  XOR31 U72215 ( .A(N3638), .B(N11284), .C(\r12190/carry [5]), .Q(N1080) );
  XOR31 U72216 ( .A(N3900), .B(N11320), .C(\r13450/carry [5]), .Q(N1110) );
  INV3 U72217 ( .A(n65781), .Q(n65758) );
  NOR21 U72218 ( .A(n66472), .B(N2103), .Q(n3364) );
  INV3 U72219 ( .A(n65607), .Q(n65602) );
  INV3 U72220 ( .A(n65584), .Q(n65577) );
  INV3 U72221 ( .A(n65606), .Q(n65603) );
  INV3 U72222 ( .A(n2358), .Q(n65444) );
  INV3 U72223 ( .A(n65611), .Q(n65609) );
  INV3 U72224 ( .A(n2060), .Q(n65440) );
  INV3 U72225 ( .A(n1890), .Q(n65442) );
  NOR31 U72226 ( .A(N1361), .B(N1300), .C(n66536), .Q(n3381) );
  NOR21 U72227 ( .A(n1691), .B(n66572), .Q(n3344) );
  NOR31 U72228 ( .A(n3649), .B(N1360), .C(n66494), .Q(n3587) );
  NAND41 U72229 ( .A(n3008), .B(n3009), .C(n3010), .D(n3011), .Q(n1696) );
  NOR21 U72230 ( .A(n1691), .B(n66572), .Q(n65549) );
  NOR21 U72231 ( .A(n1691), .B(n66572), .Q(n65550) );
  NOR31 U72232 ( .A(n3650), .B(N1903), .C(n66585), .Q(n3586) );
  NOR31 U72233 ( .A(N1905), .B(N1843), .C(N1904), .Q(n3531) );
  NOR31 U72234 ( .A(N1904), .B(N1905), .C(n66594), .Q(n3562) );
  BUF2 U72235 ( .A(n3422), .Q(n65548) );
  NOR21 U72236 ( .A(n1654), .B(state[1]), .Q(N2631) );
  BUF2 U72237 ( .A(n[5]), .Q(n65600) );
  BUF2 U72238 ( .A(\OFill[22][0] ), .Q(n65650) );
  BUF2 U72239 ( .A(\OFill[6][0] ), .Q(n65666) );
  BUF2 U72240 ( .A(\OFill[54][0] ), .Q(n65618) );
  BUF2 U72241 ( .A(\OFill[38][0] ), .Q(n65634) );
  BUF2 U72242 ( .A(\GFill[22][0] ), .Q(n65714) );
  BUF2 U72243 ( .A(\GFill[6][0] ), .Q(n65730) );
  BUF2 U72244 ( .A(\GFill[54][0] ), .Q(n65682) );
  BUF2 U72245 ( .A(\GFill[38][0] ), .Q(n65698) );
  BUF2 U72246 ( .A(\OFill[18][0] ), .Q(n65646) );
  BUF2 U72247 ( .A(\OFill[30][0] ), .Q(n65658) );
  BUF2 U72248 ( .A(\OFill[26][0] ), .Q(n65654) );
  BUF2 U72249 ( .A(\OFill[2][0] ), .Q(n65662) );
  BUF2 U72250 ( .A(\OFill[14][0] ), .Q(n65674) );
  BUF2 U72251 ( .A(\OFill[10][0] ), .Q(n65670) );
  BUF2 U72252 ( .A(\OFill[50][0] ), .Q(n65614) );
  BUF2 U72253 ( .A(\OFill[62][0] ), .Q(n65626) );
  BUF2 U72254 ( .A(\OFill[58][0] ), .Q(n65622) );
  BUF2 U72255 ( .A(\OFill[34][0] ), .Q(n65630) );
  BUF2 U72256 ( .A(\OFill[46][0] ), .Q(n65642) );
  BUF2 U72257 ( .A(\OFill[42][0] ), .Q(n65638) );
  BUF2 U72258 ( .A(\GFill[18][0] ), .Q(n65710) );
  BUF2 U72259 ( .A(\GFill[30][0] ), .Q(n65722) );
  BUF2 U72260 ( .A(\GFill[26][0] ), .Q(n65718) );
  BUF2 U72261 ( .A(\GFill[2][0] ), .Q(n65726) );
  BUF2 U72262 ( .A(\GFill[14][0] ), .Q(n65738) );
  BUF2 U72263 ( .A(\GFill[10][0] ), .Q(n65734) );
  BUF2 U72264 ( .A(\GFill[50][0] ), .Q(n65678) );
  BUF2 U72265 ( .A(\GFill[62][0] ), .Q(n65690) );
  BUF2 U72266 ( .A(\GFill[58][0] ), .Q(n65686) );
  BUF2 U72267 ( .A(\GFill[34][0] ), .Q(n65694) );
  BUF2 U72268 ( .A(\GFill[46][0] ), .Q(n65706) );
  BUF2 U72269 ( .A(\GFill[42][0] ), .Q(n65702) );
  BUF2 U72270 ( .A(n65912), .Q(n65911) );
  BUF2 U72271 ( .A(n65923), .Q(n65922) );
  BUF2 U72272 ( .A(N1130), .Q(n65538) );
  BUF2 U72273 ( .A(N1148), .Q(n65537) );
  BUF2 U72274 ( .A(N860), .Q(n65534) );
  BUF2 U72275 ( .A(n65932), .Q(n65931) );
  BUF2 U72276 ( .A(N1220), .Q(n65743) );
  BUF2 U72277 ( .A(N1082), .Q(n65912) );
  BUF2 U72278 ( .A(N1082), .Q(n65923) );
  BUF2 U72279 ( .A(N1172), .Q(n65914) );
  BUF2 U72280 ( .A(N1112), .Q(n65921) );
  BUF2 U72281 ( .A(N1184), .Q(n65913) );
  NOR21 U72282 ( .A(N2061), .B(N2060), .Q(n3618) );
  NOR21 U72283 ( .A(N1518), .B(N1517), .Q(n3614) );
  NOR20 U72284 ( .A(n66370), .B(N2061), .Q(n3525) );
  NOR20 U72285 ( .A(n66363), .B(N1518), .Q(n3523) );
  INV3 U72286 ( .A(N1517), .Q(n66363) );
  INV3 U72287 ( .A(N2060), .Q(n66370) );
  INV3 U72288 ( .A(n65437), .Q(N842) );
  BUF2 U72289 ( .A(N698), .Q(n65536) );
  BUF2 U72290 ( .A(N692), .Q(n65535) );
  BUF2 U72291 ( .A(N1016), .Q(n65933) );
  INV3 U72292 ( .A(n3470), .Q(n66369) );
  NAND20 U72293 ( .A(N2061), .B(n66370), .Q(n3470) );
  INV3 U72294 ( .A(n3466), .Q(n66362) );
  NAND20 U72295 ( .A(N1518), .B(n66363), .Q(n3466) );
  BUF2 U72296 ( .A(n65925), .Q(n65924) );
  BUF2 U72297 ( .A(n65929), .Q(n65928) );
  BUF2 U72298 ( .A(n65927), .Q(n65926) );
  BUF2 U72299 ( .A(n65935), .Q(n65934) );
  INV3 U72300 ( .A(n66109), .Q(n66114) );
  INV3 U72301 ( .A(n66098), .Q(n66103) );
  INV3 U72302 ( .A(n66092), .Q(n66097) );
  INV3 U72303 ( .A(n3377), .Q(n66477) );
  BUF2 U72304 ( .A(N1016), .Q(n65932) );
  INV3 U72305 ( .A(n65438), .Q(N1082) );
  NAND42 U72306 ( .A(N1952), .B(n66308), .C(n66314), .D(n66313), .Q(n3230) );
  NAND42 U72307 ( .A(N1409), .B(n66235), .C(n66241), .D(n66240), .Q(n3256) );
  NAND42 U72308 ( .A(n66308), .B(n66314), .C(n66313), .D(n66312), .Q(n3234) );
  NAND42 U72309 ( .A(n66235), .B(n66241), .C(n66240), .D(n66239), .Q(n3260) );
  NAND22 U72310 ( .A(n65533), .B(N11206), .Q(n3408) );
  INV0 U72311 ( .A(N11206), .Q(N1515) );
  NAND22 U72312 ( .A(n66573), .B(n3473), .Q(n3390) );
  NAND22 U72313 ( .A(n66573), .B(n3456), .Q(n3377) );
  NAND22 U72314 ( .A(n65522), .B(n66372), .Q(n3398) );
  NAND22 U72315 ( .A(N1515), .B(n65533), .Q(n3373) );
  INV6 U72316 ( .A(n65539), .Q(n65540) );
  NAND22 U72317 ( .A(n65532), .B(n66539), .Q(n3395) );
  INV3 U72318 ( .A(N1949), .Q(n66315) );
  INV3 U72319 ( .A(N1406), .Q(n66242) );
  INV6 U72320 ( .A(n65542), .Q(n65543) );
  INV6 U72321 ( .A(n65539), .Q(n65541) );
  NOR40 U72322 ( .A(n66310), .B(N1965), .C(N1967), .D(N1966), .Q(n3238) );
  INV3 U72323 ( .A(n3241), .Q(n66310) );
  NOR40 U72324 ( .A(N1971), .B(N1970), .C(N1969), .D(N1968), .Q(n3241) );
  NOR40 U72325 ( .A(n66237), .B(N1422), .C(N1424), .D(N1423), .Q(n3264) );
  INV3 U72326 ( .A(n3267), .Q(n66237) );
  NOR40 U72327 ( .A(N1428), .B(N1427), .C(N1426), .D(N1425), .Q(n3267) );
  NAND22 U72328 ( .A(n3525), .B(n3469), .Q(n3542) );
  NAND22 U72329 ( .A(n3523), .B(n3465), .Q(n3540) );
  NAND22 U72330 ( .A(n3618), .B(n3413), .Q(n3583) );
  NAND22 U72331 ( .A(n3614), .B(n3409), .Q(n3581) );
  INV3 U72332 ( .A(N1952), .Q(n66312) );
  INV3 U72333 ( .A(N1409), .Q(n66239) );
  NAND22 U72334 ( .A(n3523), .B(n3409), .Q(n3484) );
  NAND22 U72335 ( .A(n3525), .B(n3413), .Q(n3486) );
  NAND22 U72336 ( .A(n66573), .B(n3364), .Q(n3535) );
  NAND22 U72337 ( .A(n3618), .B(n3469), .Q(n3634) );
  NAND22 U72338 ( .A(n3614), .B(n3465), .Q(n3629) );
  NAND22 U72339 ( .A(n3469), .B(n66369), .Q(n3432) );
  NAND22 U72340 ( .A(n3465), .B(n66362), .Q(n3430) );
  NAND22 U72341 ( .A(n3413), .B(n66369), .Q(n3353) );
  NAND22 U72342 ( .A(n3409), .B(n66362), .Q(n3349) );
  NAND22 U72343 ( .A(n3620), .B(n3471), .Q(n3635) );
  NAND22 U72344 ( .A(n3616), .B(n3467), .Q(n3630) );
  INV3 U72345 ( .A(n65573), .Q(n65571) );
  INV3 U72346 ( .A(n65573), .Q(n65572) );
  INV3 U72347 ( .A(n65775), .Q(n65757) );
  INV3 U72348 ( .A(n65761), .Q(n65745) );
  INV3 U72349 ( .A(n65769), .Q(n65750) );
  INV3 U72350 ( .A(n65770), .Q(n65751) );
  INV3 U72351 ( .A(n65773), .Q(n65753) );
  INV3 U72352 ( .A(n65779), .Q(n65746) );
  INV3 U72353 ( .A(n65775), .Q(n65749) );
  INV3 U72354 ( .A(n65763), .Q(n65754) );
  INV3 U72355 ( .A(n65766), .Q(n65744) );
  INV3 U72356 ( .A(n65767), .Q(n65748) );
  INV3 U72357 ( .A(n65765), .Q(n65756) );
  INV3 U72358 ( .A(n65768), .Q(n65747) );
  INV3 U72359 ( .A(n65779), .Q(n65755) );
  INV3 U72360 ( .A(n65779), .Q(n65752) );
  NAND22 U72361 ( .A(n3620), .B(n3414), .Q(n3582) );
  NAND22 U72362 ( .A(n3616), .B(n3410), .Q(n3580) );
  NAND22 U72363 ( .A(n3526), .B(n3471), .Q(n3541) );
  NAND22 U72364 ( .A(n3524), .B(n3467), .Q(n3539) );
  NAND22 U72365 ( .A(n3526), .B(n3414), .Q(n3485) );
  NAND22 U72366 ( .A(n3524), .B(n3410), .Q(n3483) );
  NAND22 U72367 ( .A(n3471), .B(n66391), .Q(n3431) );
  NAND22 U72368 ( .A(n3467), .B(n66373), .Q(n3429) );
  NAND22 U72369 ( .A(n3414), .B(n66391), .Q(n3351) );
  NAND22 U72370 ( .A(n3410), .B(n66373), .Q(n3347) );
  BUF2 U72371 ( .A(n65898), .Q(n65833) );
  BUF2 U72372 ( .A(n65898), .Q(n65832) );
  BUF2 U72373 ( .A(n65898), .Q(n65834) );
  BUF2 U72374 ( .A(n65897), .Q(n65835) );
  INV3 U72375 ( .A(n3571), .Q(n66468) );
  BUF2 U72376 ( .A(n65896), .Q(n65839) );
  BUF2 U72377 ( .A(n65896), .Q(n65840) );
  BUF2 U72378 ( .A(n65896), .Q(n65838) );
  BUF2 U72379 ( .A(n65897), .Q(n65837) );
  BUF2 U72380 ( .A(n65897), .Q(n65836) );
  BUF2 U72381 ( .A(n65895), .Q(n65841) );
  BUF2 U72382 ( .A(n65895), .Q(n65842) );
  BUF2 U72383 ( .A(n65885), .Q(n65873) );
  BUF2 U72384 ( .A(n65865), .Q(n65872) );
  BUF2 U72385 ( .A(n65885), .Q(n65874) );
  BUF2 U72386 ( .A(n65892), .Q(n65850) );
  BUF2 U72387 ( .A(n65887), .Q(n65869) );
  BUF2 U72388 ( .A(n65892), .Q(n65851) );
  BUF2 U72389 ( .A(n65886), .Q(n65856) );
  BUF2 U72390 ( .A(n65849), .Q(n65855) );
  BUF2 U72391 ( .A(n65886), .Q(n65871) );
  BUF2 U72392 ( .A(n65886), .Q(n65870) );
  BUF2 U72393 ( .A(n65892), .Q(n65852) );
  BUF2 U72394 ( .A(n65891), .Q(n65854) );
  BUF2 U72395 ( .A(n65894), .Q(n65846) );
  BUF2 U72396 ( .A(n65894), .Q(n65844) );
  BUF2 U72397 ( .A(n65894), .Q(n65845) );
  BUF2 U72398 ( .A(n65893), .Q(n65847) );
  BUF2 U72399 ( .A(n65893), .Q(n65849) );
  BUF2 U72400 ( .A(n65891), .Q(n65853) );
  BUF2 U72401 ( .A(n65895), .Q(n65843) );
  BUF2 U72402 ( .A(n65892), .Q(n65858) );
  BUF2 U72403 ( .A(n65881), .Q(n65857) );
  BUF2 U72404 ( .A(n65890), .Q(n65860) );
  BUF2 U72405 ( .A(n65890), .Q(n65859) );
  BUF2 U72406 ( .A(n65889), .Q(n65863) );
  BUF2 U72407 ( .A(n65890), .Q(n65861) );
  BUF2 U72408 ( .A(n65889), .Q(n65862) );
  BUF2 U72409 ( .A(n65888), .Q(n65867) );
  BUF2 U72410 ( .A(n65887), .Q(n65868) );
  BUF2 U72411 ( .A(n65893), .Q(n65848) );
  BUF2 U72412 ( .A(n65889), .Q(n65864) );
  BUF2 U72413 ( .A(n65888), .Q(n65865) );
  BUF2 U72414 ( .A(n65888), .Q(n65866) );
  INV3 U72415 ( .A(n3489), .Q(n66473) );
  INV3 U72416 ( .A(n3358), .Q(n66395) );
  BUF2 U72417 ( .A(n65884), .Q(n65875) );
  BUF2 U72418 ( .A(n65845), .Q(n65879) );
  BUF2 U72419 ( .A(n65837), .Q(n65878) );
  BUF2 U72420 ( .A(n65866), .Q(n65876) );
  BUF2 U72421 ( .A(n65844), .Q(n65877) );
  INV3 U72422 ( .A(n3642), .Q(n66398) );
  INV3 U72423 ( .A(n3382), .Q(n66399) );
  INV3 U72424 ( .A(n66075), .Q(n66079) );
  INV3 U72425 ( .A(n66065), .Q(n66069) );
  INV3 U72426 ( .A(n3324), .Q(n66397) );
  INV3 U72427 ( .A(n3242), .Q(n66311) );
  NOR40 U72428 ( .A(N1964), .B(N1963), .C(N1962), .D(N1961), .Q(n3242) );
  INV3 U72429 ( .A(n3268), .Q(n66238) );
  NOR40 U72430 ( .A(N1421), .B(N1420), .C(N1419), .D(N1418), .Q(n3268) );
  BUF2 U72431 ( .A(n66434), .Q(n65565) );
  INV3 U72432 ( .A(n3567), .Q(n66470) );
  BUF2 U72433 ( .A(N1040), .Q(n65927) );
  BUF2 U72434 ( .A(N1046), .Q(n65925) );
  BUF2 U72435 ( .A(N1034), .Q(n65929) );
  BUF2 U72436 ( .A(N1022), .Q(n65930) );
  BUF2 U72437 ( .A(N998), .Q(n65935) );
  INV3 U72438 ( .A(N2841), .Q(n66245) );
  INV3 U72439 ( .A(N2843), .Q(n66247) );
  INV3 U72440 ( .A(N2845), .Q(n66249) );
  INV3 U72441 ( .A(N2781), .Q(n66176) );
  INV3 U72442 ( .A(N2779), .Q(n66174) );
  INV3 U72443 ( .A(N2777), .Q(n66172) );
  INV3 U72444 ( .A(N2817), .Q(n66269) );
  INV3 U72445 ( .A(N2819), .Q(n66271) );
  INV3 U72446 ( .A(N2821), .Q(n66273) );
  INV3 U72447 ( .A(N2823), .Q(n66275) );
  INV3 U72448 ( .A(N2825), .Q(n66261) );
  INV3 U72449 ( .A(N2827), .Q(n66263) );
  INV3 U72450 ( .A(N2829), .Q(n66265) );
  INV3 U72451 ( .A(N2831), .Q(n66267) );
  INV3 U72452 ( .A(N2833), .Q(n66253) );
  INV3 U72453 ( .A(N2835), .Q(n66255) );
  INV3 U72454 ( .A(N2837), .Q(n66257) );
  INV3 U72455 ( .A(N2839), .Q(n66259) );
  INV3 U72456 ( .A(N2775), .Q(n66186) );
  INV3 U72457 ( .A(N2773), .Q(n66184) );
  INV3 U72458 ( .A(N2771), .Q(n66182) );
  INV3 U72459 ( .A(N2769), .Q(n66180) );
  INV3 U72460 ( .A(N2767), .Q(n66194) );
  INV3 U72461 ( .A(N2765), .Q(n66192) );
  INV3 U72462 ( .A(N2763), .Q(n66190) );
  INV3 U72463 ( .A(N2761), .Q(n66188) );
  INV3 U72464 ( .A(N2759), .Q(n66202) );
  INV3 U72465 ( .A(N2757), .Q(n66200) );
  INV3 U72466 ( .A(N2755), .Q(n66198) );
  INV3 U72467 ( .A(N2753), .Q(n66196) );
  INV3 U72468 ( .A(N2801), .Q(n66285) );
  INV3 U72469 ( .A(N2803), .Q(n66287) );
  INV3 U72470 ( .A(N2805), .Q(n66289) );
  INV3 U72471 ( .A(N2807), .Q(n66291) );
  INV3 U72472 ( .A(N2809), .Q(n66277) );
  INV3 U72473 ( .A(N2811), .Q(n66279) );
  INV3 U72474 ( .A(N2813), .Q(n66281) );
  INV3 U72475 ( .A(N2815), .Q(n66283) );
  INV3 U72476 ( .A(N2751), .Q(n66210) );
  INV3 U72477 ( .A(N2749), .Q(n66208) );
  INV3 U72478 ( .A(N2747), .Q(n66206) );
  INV3 U72479 ( .A(N2745), .Q(n66204) );
  INV3 U72480 ( .A(N2743), .Q(n66218) );
  INV3 U72481 ( .A(N2741), .Q(n66216) );
  INV3 U72482 ( .A(N2739), .Q(n66214) );
  INV3 U72483 ( .A(N2737), .Q(n66212) );
  INV3 U72484 ( .A(N2793), .Q(n66293) );
  INV3 U72485 ( .A(N2795), .Q(n66295) );
  INV3 U72486 ( .A(N2797), .Q(n66297) );
  INV3 U72487 ( .A(N2799), .Q(n66299) );
  INV3 U72488 ( .A(N2735), .Q(n66226) );
  INV3 U72489 ( .A(N2733), .Q(n66224) );
  INV3 U72490 ( .A(N2731), .Q(n66222) );
  INV3 U72491 ( .A(N2729), .Q(n66220) );
  INV3 U72492 ( .A(N2785), .Q(n66301) );
  INV3 U72493 ( .A(N2787), .Q(n66303) );
  INV3 U72494 ( .A(N2789), .Q(n66305) );
  INV3 U72495 ( .A(N2791), .Q(n66307) );
  INV3 U72496 ( .A(N2727), .Q(n66234) );
  INV3 U72497 ( .A(N2725), .Q(n66232) );
  INV3 U72498 ( .A(N2723), .Q(n66230) );
  INV3 U72499 ( .A(N2721), .Q(n66228) );
  INV3 U72500 ( .A(N2847), .Q(n66251) );
  INV3 U72501 ( .A(N2783), .Q(n66178) );
  BUF2 U72502 ( .A(n66478), .Q(n65566) );
  NAND42 U72503 ( .A(N1952), .B(N1950), .C(n66308), .D(n66313), .Q(n3229) );
  NAND42 U72504 ( .A(N1952), .B(N1951), .C(n66308), .D(n66314), .Q(n3228) );
  NAND42 U72505 ( .A(N1409), .B(N1408), .C(n66235), .D(n66241), .Q(n3254) );
  NAND42 U72506 ( .A(N1409), .B(N1407), .C(n66235), .D(n66240), .Q(n3255) );
  NAND42 U72507 ( .A(N1951), .B(n66308), .C(n66314), .D(n66312), .Q(n3232) );
  NAND42 U72508 ( .A(N1951), .B(N1950), .C(n66308), .D(n66312), .Q(n3231) );
  NAND42 U72509 ( .A(N1408), .B(N1407), .C(n66235), .D(n66239), .Q(n3257) );
  NAND42 U72510 ( .A(N1408), .B(n66235), .C(n66241), .D(n66239), .Q(n3258) );
  NAND42 U72511 ( .A(N1950), .B(n66308), .C(n66313), .D(n66312), .Q(n3233) );
  NAND42 U72512 ( .A(N1407), .B(n66235), .C(n66240), .D(n66239), .Q(n3259) );
  NAND42 U72513 ( .A(N1952), .B(N1951), .C(N1950), .D(n66308), .Q(n3220) );
  NAND42 U72514 ( .A(N1409), .B(N1408), .C(N1407), .D(n66235), .Q(n3246) );
  XNR21 U72515 ( .A(n65602), .B(n65578), .Q(N3899) );
  NAND33 U72516 ( .A(N1947), .B(n66316), .C(N1949), .Q(n3222) );
  NAND33 U72517 ( .A(N1404), .B(n66243), .C(N1406), .Q(n3248) );
  NAND33 U72518 ( .A(N1948), .B(N1947), .C(N1949), .Q(n3219) );
  NAND33 U72519 ( .A(N1405), .B(N1404), .C(N1406), .Q(n3245) );
  NAND33 U72520 ( .A(N1947), .B(n66315), .C(N1948), .Q(n3224) );
  NAND33 U72521 ( .A(N1404), .B(n66242), .C(N1405), .Q(n3250) );
  NAND33 U72522 ( .A(n66316), .B(n66315), .C(N1947), .Q(n3226) );
  NAND33 U72523 ( .A(n66243), .B(n66242), .C(N1404), .Q(n3252) );
  NOR22 U72524 ( .A(n3639), .B(n3571), .Q(n3386) );
  NAND22 U72525 ( .A(N2058), .B(n65518), .Q(n3354) );
  NOR21 U72526 ( .A(n66487), .B(n66471), .Q(n3421) );
  NOR21 U72527 ( .A(n66472), .B(n66569), .Q(n3473) );
  NOR21 U72528 ( .A(n66569), .B(n65576), .Q(n3456) );
  INV3 U72529 ( .A(N2058), .Q(n66372) );
  NOR21 U72530 ( .A(n3571), .B(n66484), .Q(n3336) );
  INV3 U72531 ( .A(n3561), .Q(n66484) );
  NAND22 U72532 ( .A(n3473), .B(n3563), .Q(n3341) );
  INV3 U72533 ( .A(n66110), .Q(N1041) );
  INV3 U72534 ( .A(n66088), .Q(N1047) );
  INV3 U72535 ( .A(n66084), .Q(N1035) );
  INV3 U72536 ( .A(n66115), .Q(N1017) );
  INV3 U72537 ( .A(n66099), .Q(N1023) );
  INV3 U72538 ( .A(n66093), .Q(N999) );
  NOR21 U72539 ( .A(n3619), .B(N2059), .Q(n3469) );
  NOR21 U72540 ( .A(n3615), .B(N1516), .Q(n3465) );
  NOR21 U72541 ( .A(n65573), .B(N1560), .Q(n3358) );
  NAND22 U72542 ( .A(n3456), .B(n3563), .Q(n3331) );
  NAND22 U72543 ( .A(n66398), .B(n3561), .Q(n3324) );
  INV3 U72544 ( .A(N1946), .Q(n65542) );
  INV3 U72545 ( .A(N1403), .Q(n65539) );
  NOR40 U72546 ( .A(n3243), .B(N1955), .C(N1957), .D(N1956), .Q(n3236) );
  NAND22 U72547 ( .A(n3244), .B(n66478), .Q(n3243) );
  NOR21 U72548 ( .A(N1954), .B(N1953), .Q(n3244) );
  NOR40 U72549 ( .A(n3269), .B(N1412), .C(N1414), .D(N1413), .Q(n3262) );
  NAND22 U72550 ( .A(n3270), .B(n66434), .Q(n3269) );
  NOR21 U72551 ( .A(N1411), .B(N1410), .Q(n3270) );
  INV3 U72552 ( .A(n3235), .Q(n66308) );
  NAND41 U72553 ( .A(n3236), .B(n3237), .C(n3238), .D(n3239), .Q(n3235) );
  NOR40 U72554 ( .A(n66309), .B(N1972), .C(N1974), .D(N1973), .Q(n3239) );
  NOR40 U72555 ( .A(n66311), .B(N1958), .C(N1960), .D(N1959), .Q(n3237) );
  INV3 U72556 ( .A(n3261), .Q(n66235) );
  NAND41 U72557 ( .A(n3262), .B(n3263), .C(n3264), .D(n3265), .Q(n3261) );
  NOR40 U72558 ( .A(n66236), .B(N1429), .C(N1431), .D(N1430), .Q(n3265) );
  NOR40 U72559 ( .A(n66238), .B(N1415), .C(N1417), .D(N1416), .Q(n3263) );
  NOR40 U72560 ( .A(N1315), .B(N1314), .C(N1313), .D(N1312), .Q(n66866) );
  NOR40 U72561 ( .A(N1305), .B(N1304), .C(N1303), .D(N1330), .Q(n66861) );
  NOR40 U72562 ( .A(N1329), .B(N1328), .C(N1327), .D(N1326), .Q(n66862) );
  NOR40 U72563 ( .A(N1858), .B(N1857), .C(N1856), .D(N1855), .Q(n66880) );
  NOR40 U72564 ( .A(N1848), .B(N1847), .C(N1846), .D(N1873), .Q(n66875) );
  NOR40 U72565 ( .A(N1872), .B(N1871), .C(N1870), .D(N1869), .Q(n66876) );
  NAND22 U72566 ( .A(N1526), .B(n65532), .Q(n3348) );
  NAND22 U72567 ( .A(n65451), .B(n65522), .Q(n3374) );
  NAND22 U72568 ( .A(N1910), .B(n3279), .Q(n3271) );
  NOR40 U72569 ( .A(N1309), .B(N1308), .C(N1307), .D(N1306), .Q(n66860) );
  NOR40 U72570 ( .A(N1852), .B(N1851), .C(N1850), .D(N1849), .Q(n66874) );
  NAND22 U72571 ( .A(n3279), .B(n66645), .Q(n3280) );
  INV3 U72572 ( .A(N1910), .Q(n66645) );
  NOR21 U72573 ( .A(n65576), .B(N2103), .Q(n3489) );
  NOR21 U72574 ( .A(n3639), .B(n3642), .Q(n3382) );
  NOR40 U72575 ( .A(n66504), .B(N1316), .C(N1318), .D(N1317), .Q(n66865) );
  INV3 U72576 ( .A(n66864), .Q(n66504) );
  NOR40 U72577 ( .A(N1322), .B(N1321), .C(N1320), .D(N1319), .Q(n66864) );
  NOR40 U72578 ( .A(n66593), .B(N1859), .C(N1861), .D(N1860), .Q(n66879) );
  INV3 U72579 ( .A(n66878), .Q(n66593) );
  NOR40 U72580 ( .A(N1865), .B(N1864), .C(N1863), .D(N1862), .Q(n66878) );
  NAND22 U72581 ( .A(n66469), .B(N1560), .Q(n3571) );
  XOR21 U72582 ( .A(m[2]), .B(n66651), .Q(N5356) );
  NAND22 U72583 ( .A(n65577), .B(n65604), .Q(n66651) );
  XOR21 U72584 ( .A(m[2]), .B(n66650), .Q(N3086) );
  NAND22 U72585 ( .A(n65577), .B(m[1]), .Q(n66650) );
  INV3 U72586 ( .A(N4602), .Q(n66564) );
  INV3 U72587 ( .A(N1948), .Q(n66316) );
  INV3 U72588 ( .A(N1405), .Q(n66243) );
  NAND22 U72589 ( .A(N1560), .B(n65571), .Q(n3642) );
  INV3 U72590 ( .A(N1951), .Q(n66313) );
  INV3 U72591 ( .A(N1408), .Q(n66240) );
  INV3 U72592 ( .A(n66127), .Q(N1029) );
  INV3 U72593 ( .A(n66135), .Q(N1011) );
  INV3 U72594 ( .A(n66139), .Q(N1005) );
  INV3 U72595 ( .A(n66151), .Q(N993) );
  INV3 U72596 ( .A(n66159), .Q(N981) );
  INV3 U72597 ( .A(n66155), .Q(N987) );
  INV3 U72598 ( .A(n66131), .Q(N741) );
  INV3 U72599 ( .A(n66143), .Q(N723) );
  INV3 U72600 ( .A(n66147), .Q(N717) );
  INV3 U72601 ( .A(n66163), .Q(N705) );
  INV3 U72602 ( .A(N1950), .Q(n66314) );
  INV3 U72603 ( .A(N1407), .Q(n66241) );
  NOR21 U72604 ( .A(n66480), .B(n3278), .Q(n3273) );
  INV3 U72605 ( .A(N1367), .Q(n66480) );
  NOR21 U72606 ( .A(n3278), .B(N1367), .Q(n3282) );
  XNR21 U72607 ( .A(m[2]), .B(n65602), .Q(N6300) );
  XNR21 U72608 ( .A(n65609), .B(n65602), .Q(N5511) );
  XNR21 U72609 ( .A(m[2]), .B(n65602), .Q(N5338) );
  XNR21 U72610 ( .A(n65609), .B(n65602), .Q(N3241) );
  XNR21 U72611 ( .A(n65609), .B(n65602), .Q(N3068) );
  XNR21 U72612 ( .A(m[2]), .B(n65603), .Q(N6437) );
  XNR21 U72613 ( .A(m[2]), .B(n65603), .Q(N6576) );
  XNR21 U72614 ( .A(n65609), .B(n65603), .Q(N7266) );
  XNR21 U72615 ( .A(m[2]), .B(n65603), .Q(N4167) );
  XNR21 U72616 ( .A(m[2]), .B(n65603), .Q(N4306) );
  XNR21 U72617 ( .A(n65609), .B(n65603), .Q(N4996) );
  XNR21 U72618 ( .A(m[2]), .B(n65603), .Q(N7013) );
  XNR21 U72619 ( .A(m[2]), .B(n65603), .Q(N4743) );
  NOR21 U72620 ( .A(n66371), .B(n3619), .Q(n3413) );
  INV3 U72621 ( .A(N2059), .Q(n66371) );
  NOR21 U72622 ( .A(n66364), .B(n3615), .Q(n3409) );
  INV3 U72623 ( .A(N1516), .Q(n66364) );
  NOR21 U72624 ( .A(n3621), .B(N2070), .Q(n3471) );
  NOR21 U72625 ( .A(n66487), .B(n3642), .Q(n3504) );
  NOR21 U72626 ( .A(n3617), .B(N1527), .Q(n3467) );
  BUF2 U72627 ( .A(N4855), .Q(n65555) );
  XNR21 U72628 ( .A(n65609), .B(n3180), .Q(N4855) );
  NAND22 U72629 ( .A(n65604), .B(n65578), .Q(n3180) );
  NOR21 U72630 ( .A(n66644), .B(n3621), .Q(n3414) );
  INV3 U72631 ( .A(N2070), .Q(n66644) );
  NOR21 U72632 ( .A(n66479), .B(n3617), .Q(n3410) );
  INV3 U72633 ( .A(N1527), .Q(n66479) );
  NOR31 U72634 ( .A(N1323), .B(N1325), .C(N1324), .Q(n66863) );
  NOR31 U72635 ( .A(N1866), .B(N1868), .C(N1867), .Q(n66877) );
  INV3 U72636 ( .A(n3383), .Q(n66527) );
  INV3 U72637 ( .A(n3641), .Q(n66588) );
  NOR21 U72638 ( .A(n3639), .B(n66471), .Q(n3567) );
  NOR21 U72639 ( .A(n3639), .B(n66395), .Q(n3529) );
  BUF6 U72640 ( .A(n66568), .Q(n65568) );
  BUF6 U72641 ( .A(n66568), .Q(n65567) );
  BUF2 U72642 ( .A(n65949), .Q(n65953) );
  BUF2 U72643 ( .A(n65939), .Q(n65943) );
  BUF2 U72644 ( .A(n65948), .Q(n65952) );
  BUF2 U72645 ( .A(n65938), .Q(n65942) );
  BUF2 U72646 ( .A(n65940), .Q(n65944) );
  BUF2 U72647 ( .A(n65950), .Q(n65954) );
  AOI211 U72648 ( .A(n65604), .B(n65577), .C(n65610), .Q(n66825) );
  AOI211 U72649 ( .A(n65604), .B(n65577), .C(n65610), .Q(n66740) );
  NOR21 U72650 ( .A(n3640), .B(n66473), .Q(n3530) );
  NAND22 U72651 ( .A(n65577), .B(N4857), .Q(n66678) );
  NAND22 U72652 ( .A(n65577), .B(N3395), .Q(n66657) );
  NAND22 U72653 ( .A(n65577), .B(N3359), .Q(n66655) );
  NAND22 U72654 ( .A(n65579), .B(N3222), .Q(n66654) );
  NAND22 U72655 ( .A(n65578), .B(N3049), .Q(n66652) );
  NAND22 U72656 ( .A(n65577), .B(N4718), .Q(n66674) );
  NAND22 U72657 ( .A(n65577), .B(N4605), .Q(n66673) );
  NAND22 U72658 ( .A(n65577), .B(N4581), .Q(n66671) );
  NAND22 U72659 ( .A(n65577), .B(N4468), .Q(n66670) );
  INV3 U72660 ( .A(n3594), .Q(n66590) );
  NAND31 U72661 ( .A(n65757), .B(n65835), .C(n65915), .Q(n66842) );
  BUF2 U72662 ( .A(n65453), .Q(n65533) );
  BUF2 U72663 ( .A(n65514), .Q(n65516) );
  BUF2 U72664 ( .A(n65531), .Q(n65530) );
  BUF2 U72665 ( .A(n65419), .Q(n65512) );
  BUF2 U72666 ( .A(n65419), .Q(n65511) );
  BUF2 U72667 ( .A(n65453), .Q(n65524) );
  BUF2 U72668 ( .A(n65524), .Q(n65528) );
  BUF2 U72669 ( .A(n65532), .Q(n65529) );
  BUF2 U72670 ( .A(n65419), .Q(n65513) );
  BUF2 U72671 ( .A(n65520), .Q(n65519) );
  BUF2 U72672 ( .A(n65512), .Q(n65518) );
  BUF2 U72673 ( .A(n65419), .Q(n65510) );
  BUF2 U72674 ( .A(n65517), .Q(n65515) );
  BUF2 U72675 ( .A(n65511), .Q(n65514) );
  BUF2 U72676 ( .A(n65453), .Q(n65525) );
  BUF2 U72677 ( .A(n65453), .Q(n65526) );
  BUF2 U72678 ( .A(n65453), .Q(n65523) );
  BUF2 U72679 ( .A(n65518), .Q(n65521) );
  BUF2 U72680 ( .A(n65510), .Q(n65520) );
  BUF2 U72681 ( .A(n65453), .Q(n65527) );
  BUF2 U72682 ( .A(n65513), .Q(n65517) );
  BUF2 U72683 ( .A(n65420), .Q(n65531) );
  BUF2 U72684 ( .A(n65453), .Q(n65532) );
  INV3 U72685 ( .A(n65576), .Q(n65575) );
  INV3 U72686 ( .A(n65576), .Q(n65574) );
  BUF2 U72687 ( .A(n65512), .Q(n65522) );
  BUF2 U72688 ( .A(n65883), .Q(n65881) );
  BUF2 U72689 ( .A(n65883), .Q(n65880) );
  NOR21 U72690 ( .A(n66392), .B(N2072), .Q(n3526) );
  NOR21 U72691 ( .A(n66374), .B(N1529), .Q(n3524) );
  NOR21 U72692 ( .A(N2072), .B(N2071), .Q(n3620) );
  NOR21 U72693 ( .A(N1529), .B(N1528), .Q(n3616) );
  INV3 U72694 ( .A(N2103), .Q(n66569) );
  INV3 U72695 ( .A(n3494), .Q(n66471) );
  NOR21 U72696 ( .A(N1311), .B(N1310), .Q(n66868) );
  NOR21 U72697 ( .A(N1854), .B(N1853), .Q(n66882) );
  BUF2 U72698 ( .A(n65941), .Q(n65945) );
  BUF2 U72699 ( .A(n65951), .Q(n65955) );
  INV3 U72700 ( .A(n3563), .Q(n66574) );
  NAND22 U72701 ( .A(n65578), .B(n65604), .Q(n66648) );
  NAND22 U72702 ( .A(n65577), .B(n65602), .Q(n66661) );
  INV3 U72703 ( .A(N1526), .Q(n66539) );
  INV3 U72704 ( .A(n66064), .Q(n66070) );
  INV3 U72705 ( .A(n66074), .Q(n66080) );
  BUF2 U72706 ( .A(n65774), .Q(n65773) );
  BUF2 U72707 ( .A(n65775), .Q(n65771) );
  BUF2 U72708 ( .A(n65775), .Q(n65770) );
  BUF2 U72709 ( .A(n65776), .Q(n65766) );
  BUF2 U72710 ( .A(n65777), .Q(n65765) );
  BUF2 U72711 ( .A(n65761), .Q(n65772) );
  BUF2 U72712 ( .A(n65775), .Q(n65769) );
  BUF2 U72713 ( .A(n65776), .Q(n65767) );
  BUF2 U72714 ( .A(n65776), .Q(n65768) );
  BUF2 U72715 ( .A(n65777), .Q(n65764) );
  BUF2 U72716 ( .A(n65777), .Q(n65763) );
  BUF2 U72717 ( .A(n65778), .Q(n65762) );
  BUF2 U72718 ( .A(n65778), .Q(n65760) );
  BUF2 U72719 ( .A(n65778), .Q(n65761) );
  BUF2 U72720 ( .A(n65761), .Q(n65759) );
  INV3 U72721 ( .A(N2071), .Q(n66392) );
  INV3 U72722 ( .A(N1528), .Q(n66374) );
  INV3 U72723 ( .A(n65552), .Q(n66530) );
  BUF2 U72724 ( .A(n65883), .Q(n65882) );
  INV3 U72725 ( .A(n3218), .Q(n66478) );
  INV3 U72726 ( .A(n3640), .Q(n66573) );
  INV3 U72727 ( .A(n3217), .Q(n66434) );
  INV3 U72728 ( .A(n3287), .Q(n65573) );
  INV3 U72729 ( .A(n3472), .Q(n66391) );
  NAND22 U72730 ( .A(N2072), .B(n66392), .Q(n3472) );
  INV3 U72731 ( .A(n3468), .Q(n66373) );
  NAND22 U72732 ( .A(N1529), .B(n66374), .Q(n3468) );
  INV3 U72733 ( .A(n3461), .Q(n66488) );
  INV3 U72734 ( .A(n3438), .Q(n66474) );
  INV3 U72735 ( .A(n65591), .Q(n65589) );
  INV3 U72736 ( .A(n65591), .Q(n65588) );
  INV3 U72737 ( .A(n65591), .Q(n65587) );
  INV3 U72738 ( .A(n65590), .Q(n65586) );
  BUF2 U72739 ( .A(n66393), .Q(n65564) );
  BUF2 U72740 ( .A(n66382), .Q(n65563) );
  BUF2 U72741 ( .A(n66381), .Q(n65562) );
  BUF2 U72742 ( .A(n66377), .Q(n65558) );
  BUF2 U72743 ( .A(n66378), .Q(n65559) );
  BUF2 U72744 ( .A(n66375), .Q(n65556) );
  BUF2 U72745 ( .A(n66379), .Q(n65560) );
  BUF2 U72746 ( .A(n66376), .Q(n65557) );
  INV3 U72747 ( .A(n3360), .Q(n66396) );
  INV3 U72748 ( .A(n3682), .Q(n66335) );
  INV3 U72749 ( .A(n3602), .Q(n66351) );
  INV3 U72750 ( .A(n3628), .Q(n66340) );
  INV3 U72751 ( .A(n3646), .Q(n66338) );
  BUF2 U72752 ( .A(n65900), .Q(n65896) );
  BUF2 U72753 ( .A(n65905), .Q(n65885) );
  BUF2 U72754 ( .A(n65902), .Q(n65892) );
  BUF2 U72755 ( .A(n65906), .Q(n65884) );
  BUF2 U72756 ( .A(n65904), .Q(n65887) );
  BUF2 U72757 ( .A(n65904), .Q(n65886) );
  BUF2 U72758 ( .A(n65901), .Q(n65894) );
  BUF2 U72759 ( .A(n65902), .Q(n65893) );
  BUF2 U72760 ( .A(n65894), .Q(n65891) );
  BUF2 U72761 ( .A(n65900), .Q(n65897) );
  BUF2 U72762 ( .A(n65848), .Q(n65890) );
  BUF2 U72763 ( .A(n65901), .Q(n65895) );
  BUF2 U72764 ( .A(n65899), .Q(n65898) );
  BUF2 U72765 ( .A(n65903), .Q(n65889) );
  BUF2 U72766 ( .A(n65903), .Q(n65888) );
  BUF2 U72767 ( .A(n66568), .Q(n65569) );
  INV3 U72768 ( .A(N2840), .Q(n66244) );
  INV3 U72769 ( .A(N2842), .Q(n66246) );
  INV3 U72770 ( .A(N2844), .Q(n66248) );
  INV3 U72771 ( .A(N2846), .Q(n66250) );
  INV3 U72772 ( .A(N2782), .Q(n66177) );
  INV3 U72773 ( .A(N2780), .Q(n66175) );
  INV3 U72774 ( .A(N2778), .Q(n66173) );
  INV3 U72775 ( .A(N2776), .Q(n66171) );
  INV3 U72776 ( .A(n3211), .Q(n66430) );
  AOI221 U72777 ( .A(N1844), .B(n65566), .C(N1301), .D(n65565), .Q(n3211) );
  INV3 U72778 ( .A(n3210), .Q(n66429) );
  AOI221 U72779 ( .A(N1845), .B(n66478), .C(N1302), .D(n66434), .Q(n3210) );
  INV3 U72780 ( .A(n3201), .Q(n66420) );
  AOI221 U72781 ( .A(N1854), .B(n65566), .C(N1311), .D(n65565), .Q(n3201) );
  INV3 U72782 ( .A(n3189), .Q(n66408) );
  AOI221 U72783 ( .A(N1866), .B(n66478), .C(N1323), .D(n66434), .Q(n3189) );
  INV3 U72784 ( .A(n3187), .Q(n66406) );
  AOI221 U72785 ( .A(N1868), .B(n65566), .C(N1325), .D(n66434), .Q(n3187) );
  INV3 U72786 ( .A(n3188), .Q(n66407) );
  AOI221 U72787 ( .A(N1867), .B(n66478), .C(N1324), .D(n66434), .Q(n3188) );
  INV3 U72788 ( .A(n3202), .Q(n66421) );
  AOI221 U72789 ( .A(N1853), .B(n66478), .C(N1310), .D(n66434), .Q(n3202) );
  INV3 U72790 ( .A(n3185), .Q(n66404) );
  AOI221 U72791 ( .A(N1870), .B(n65566), .C(N1327), .D(n65565), .Q(n3185) );
  INV3 U72792 ( .A(n3192), .Q(n66411) );
  AOI221 U72793 ( .A(N1863), .B(n66478), .C(N1320), .D(n66434), .Q(n3192) );
  INV3 U72794 ( .A(n3194), .Q(n66413) );
  AOI221 U72795 ( .A(N1861), .B(n65566), .C(N1318), .D(n65565), .Q(n3194) );
  INV3 U72796 ( .A(n3199), .Q(n66418) );
  AOI221 U72797 ( .A(N1856), .B(n66478), .C(N1313), .D(n65565), .Q(n3199) );
  INV3 U72798 ( .A(n3205), .Q(n66424) );
  AOI221 U72799 ( .A(N1850), .B(n65566), .C(N1307), .D(n66434), .Q(n3205) );
  BUF2 U72800 ( .A(n66380), .Q(n65561) );
  INV3 U72801 ( .A(n3182), .Q(n66401) );
  AOI221 U72802 ( .A(N1873), .B(n65566), .C(N1330), .D(n66434), .Q(n3182) );
  INV3 U72803 ( .A(n3184), .Q(n66403) );
  AOI221 U72804 ( .A(N1871), .B(n65566), .C(N1328), .D(n65565), .Q(n3184) );
  INV3 U72805 ( .A(n3186), .Q(n66405) );
  AOI221 U72806 ( .A(N1869), .B(n66478), .C(N1326), .D(n66434), .Q(n3186) );
  INV3 U72807 ( .A(n3191), .Q(n66410) );
  AOI221 U72808 ( .A(N1864), .B(n65566), .C(N1321), .D(n65565), .Q(n3191) );
  INV3 U72809 ( .A(n3193), .Q(n66412) );
  AOI221 U72810 ( .A(N1862), .B(n66478), .C(N1319), .D(n66434), .Q(n3193) );
  INV3 U72811 ( .A(n3195), .Q(n66414) );
  AOI221 U72812 ( .A(N1860), .B(n65566), .C(N1317), .D(n65565), .Q(n3195) );
  INV3 U72813 ( .A(n3196), .Q(n66415) );
  AOI221 U72814 ( .A(N1859), .B(n66478), .C(N1316), .D(n65565), .Q(n3196) );
  INV3 U72815 ( .A(n3198), .Q(n66417) );
  AOI221 U72816 ( .A(N1857), .B(n65566), .C(N1314), .D(n66434), .Q(n3198) );
  INV3 U72817 ( .A(n3200), .Q(n66419) );
  AOI221 U72818 ( .A(N1855), .B(n66478), .C(N1312), .D(n65565), .Q(n3200) );
  INV3 U72819 ( .A(n3204), .Q(n66423) );
  AOI221 U72820 ( .A(N1851), .B(n65566), .C(N1308), .D(n66434), .Q(n3204) );
  INV3 U72821 ( .A(n3206), .Q(n66425) );
  AOI221 U72822 ( .A(N1849), .B(n66478), .C(N1306), .D(n66434), .Q(n3206) );
  INV3 U72823 ( .A(n3208), .Q(n66427) );
  AOI221 U72824 ( .A(N1847), .B(n65566), .C(N1304), .D(n66434), .Q(n3208) );
  INV3 U72825 ( .A(n3183), .Q(n66402) );
  AOI221 U72826 ( .A(N1872), .B(n66478), .C(N1329), .D(n66434), .Q(n3183) );
  INV3 U72827 ( .A(n3190), .Q(n66409) );
  AOI221 U72828 ( .A(N1865), .B(n65566), .C(N1322), .D(n65565), .Q(n3190) );
  INV3 U72829 ( .A(n3197), .Q(n66416) );
  AOI221 U72830 ( .A(N1858), .B(n66478), .C(N1315), .D(n66434), .Q(n3197) );
  INV3 U72831 ( .A(n3203), .Q(n66422) );
  AOI221 U72832 ( .A(N1852), .B(n66478), .C(N1309), .D(n66434), .Q(n3203) );
  INV3 U72833 ( .A(n3207), .Q(n66426) );
  AOI221 U72834 ( .A(N1848), .B(n66478), .C(N1305), .D(n66434), .Q(n3207) );
  INV3 U72835 ( .A(N2816), .Q(n66268) );
  INV3 U72836 ( .A(N2818), .Q(n66270) );
  INV3 U72837 ( .A(N2820), .Q(n66272) );
  INV3 U72838 ( .A(N2822), .Q(n66274) );
  INV3 U72839 ( .A(N2824), .Q(n66260) );
  INV3 U72840 ( .A(N2826), .Q(n66262) );
  INV3 U72841 ( .A(N2828), .Q(n66264) );
  INV3 U72842 ( .A(N2830), .Q(n66266) );
  INV3 U72843 ( .A(N2832), .Q(n66252) );
  INV3 U72844 ( .A(N2834), .Q(n66254) );
  INV3 U72845 ( .A(N2836), .Q(n66256) );
  INV3 U72846 ( .A(N2838), .Q(n66258) );
  INV3 U72847 ( .A(N2774), .Q(n66185) );
  INV3 U72848 ( .A(N2772), .Q(n66183) );
  INV3 U72849 ( .A(N2770), .Q(n66181) );
  INV3 U72850 ( .A(N2768), .Q(n66179) );
  INV3 U72851 ( .A(N2766), .Q(n66193) );
  INV3 U72852 ( .A(N2764), .Q(n66191) );
  INV3 U72853 ( .A(N2762), .Q(n66189) );
  INV3 U72854 ( .A(N2760), .Q(n66187) );
  INV3 U72855 ( .A(N2758), .Q(n66201) );
  INV3 U72856 ( .A(N2756), .Q(n66199) );
  INV3 U72857 ( .A(N2754), .Q(n66197) );
  INV3 U72858 ( .A(N2752), .Q(n66195) );
  INV3 U72859 ( .A(N2800), .Q(n66284) );
  INV3 U72860 ( .A(N2802), .Q(n66286) );
  INV3 U72861 ( .A(N2804), .Q(n66288) );
  INV3 U72862 ( .A(N2806), .Q(n66290) );
  INV3 U72863 ( .A(N2808), .Q(n66276) );
  INV3 U72864 ( .A(N2810), .Q(n66278) );
  INV3 U72865 ( .A(N2812), .Q(n66280) );
  INV3 U72866 ( .A(N2814), .Q(n66282) );
  INV3 U72867 ( .A(N2750), .Q(n66209) );
  INV3 U72868 ( .A(N2748), .Q(n66207) );
  INV3 U72869 ( .A(N2746), .Q(n66205) );
  INV3 U72870 ( .A(N2744), .Q(n66203) );
  INV3 U72871 ( .A(N2742), .Q(n66217) );
  INV3 U72872 ( .A(N2740), .Q(n66215) );
  INV3 U72873 ( .A(N2738), .Q(n66213) );
  INV3 U72874 ( .A(N2736), .Q(n66211) );
  INV3 U72875 ( .A(N2792), .Q(n66292) );
  INV3 U72876 ( .A(N2794), .Q(n66294) );
  INV3 U72877 ( .A(N2796), .Q(n66296) );
  INV3 U72878 ( .A(N2798), .Q(n66298) );
  INV3 U72879 ( .A(N2734), .Q(n66225) );
  INV3 U72880 ( .A(N2732), .Q(n66223) );
  INV3 U72881 ( .A(N2730), .Q(n66221) );
  INV3 U72882 ( .A(N2728), .Q(n66219) );
  INV3 U72883 ( .A(N2784), .Q(n66300) );
  INV3 U72884 ( .A(N2786), .Q(n66302) );
  INV3 U72885 ( .A(N2788), .Q(n66304) );
  INV3 U72886 ( .A(N2790), .Q(n66306) );
  INV3 U72887 ( .A(N2726), .Q(n66233) );
  INV3 U72888 ( .A(N2724), .Q(n66231) );
  INV3 U72889 ( .A(N2722), .Q(n66229) );
  INV3 U72890 ( .A(N2720), .Q(n66227) );
  INV3 U72891 ( .A(n3209), .Q(n66428) );
  AOI221 U72892 ( .A(N1846), .B(n66478), .C(N1303), .D(n66434), .Q(n3209) );
  INV3 U72893 ( .A(N2674), .Q(n66359) );
  AOI2111 U72894 ( .A(n3386), .B(n3383), .C(n3387), .D(n3388), .Q(n3385) );
  INV3 U72895 ( .A(N2668), .Q(n66347) );
  AOI2111 U72896 ( .A(n65552), .B(n3386), .C(n3440), .D(n3441), .Q(n3439) );
  INV3 U72897 ( .A(N2634), .Q(n66336) );
  AOI2111 U72898 ( .A(n65552), .B(n3421), .C(n3658), .D(n3659), .Q(n3657) );
  NOR40 U72899 ( .A(n2315), .B(n2273), .C(n1696), .D(n66467), .Q(n1685) );
  AOI311 U72900 ( .A(n66317), .B(n1728), .C(n1729), .D(n66467), .Q(n1727) );
  INV3 U72901 ( .A(n2244), .Q(n66317) );
  NOR31 U72902 ( .A(n2102), .B(n2230), .C(n2145), .Q(n1728) );
  NOR40 U72903 ( .A(n1730), .B(n1731), .C(n1803), .D(n1761), .Q(n1729) );
  XNR21 U72904 ( .A(n65609), .B(n65607), .Q(N4728) );
  XNR21 U72905 ( .A(n65583), .B(n65602), .Q(N2913) );
  NOR32 U72906 ( .A(n66537), .B(n66531), .C(n66536), .Q(n3383) );
  XOR21 U72907 ( .A(n65610), .B(n3179), .Q(N4603) );
  NAND22 U72908 ( .A(N4602), .B(n65581), .Q(n3179) );
  INV3 U72909 ( .A(N1331), .Q(n66482) );
  NAND41 U72910 ( .A(n66863), .B(n66862), .C(n66861), .D(n66860), .Q(n66870)
         );
  NAND41 U72911 ( .A(n66868), .B(n66867), .C(n66866), .D(n66865), .Q(n66869)
         );
  NOR31 U72912 ( .A(n66526), .B(n3649), .C(n66494), .Q(n3561) );
  XOR21 U72913 ( .A(n66537), .B(n66536), .Q(N1301) );
  XOR21 U72914 ( .A(n66594), .B(n66596), .Q(N1844) );
  NAND22 U72915 ( .A(n65742), .B(N11206), .Q(n3396) );
  NAND33 U72916 ( .A(N1843), .B(n66316), .C(N1949), .Q(n3223) );
  NAND33 U72917 ( .A(N1948), .B(N1843), .C(N1949), .Q(n3221) );
  NAND33 U72918 ( .A(N1405), .B(n65546), .C(N1406), .Q(n3247) );
  NAND33 U72919 ( .A(n65546), .B(n66243), .C(N1406), .Q(n3249) );
  NAND33 U72920 ( .A(N1843), .B(n66315), .C(N1948), .Q(n3225) );
  NAND33 U72921 ( .A(n65546), .B(n66242), .C(N1405), .Q(n3251) );
  XOR21 U72922 ( .A(\sub_126_S2_2/carry [2]), .B(n66531), .Q(N1302) );
  XOR21 U72923 ( .A(\sub_157_S2_2/carry [2]), .B(n66597), .Q(N1845) );
  NAND33 U72924 ( .A(n66316), .B(n66315), .C(n65545), .Q(n3227) );
  NAND33 U72925 ( .A(n66243), .B(n66242), .C(N1300), .Q(n3253) );
  INV3 U72926 ( .A(N1874), .Q(n66570) );
  NAND41 U72927 ( .A(n66877), .B(n66876), .C(n66875), .D(n66874), .Q(n66884)
         );
  NAND41 U72928 ( .A(n66882), .B(n66881), .C(n66880), .D(n66879), .Q(n66883)
         );
  XOR21 U72929 ( .A(\sub_126_S2_2/carry [11]), .B(n66518), .Q(N1311) );
  XOR21 U72930 ( .A(\sub_157_S2_2/carry [11]), .B(n66607), .Q(N1854) );
  XOR21 U72931 ( .A(\sub_126_S2_2/carry [23]), .B(n66503), .Q(N1323) );
  XOR21 U72932 ( .A(\sub_126_S2_2/carry [25]), .B(n66500), .Q(N1325) );
  XOR21 U72933 ( .A(\sub_157_S2_2/carry [23]), .B(n66621), .Q(N1866) );
  NOR31 U72934 ( .A(n66598), .B(n3650), .C(n66585), .Q(n3563) );
  XOR21 U72935 ( .A(\sub_126_S2_2/carry [10]), .B(n66519), .Q(N1310) );
  XOR21 U72936 ( .A(\sub_126_S2_2/carry [24]), .B(n66501), .Q(N1324) );
  XOR21 U72937 ( .A(\sub_157_S2_2/carry [25]), .B(n66623), .Q(N1868) );
  XOR21 U72938 ( .A(\sub_157_S2_2/carry [10]), .B(n66605), .Q(N1853) );
  XOR21 U72939 ( .A(\sub_157_S2_2/carry [24]), .B(n66622), .Q(N1867) );
  XOR21 U72940 ( .A(\sub_126_S2_2/carry [20]), .B(n66507), .Q(N1320) );
  XOR21 U72941 ( .A(\sub_126_S2_2/carry [13]), .B(n66516), .Q(N1313) );
  XOR21 U72942 ( .A(\sub_126_S2_2/carry [18]), .B(n66509), .Q(N1318) );
  XOR21 U72943 ( .A(\sub_126_S2_2/carry [27]), .B(n66498), .Q(N1327) );
  XOR21 U72944 ( .A(\sub_126_S2_2/carry [7]), .B(n66522), .Q(N1307) );
  XOR21 U72945 ( .A(\sub_126_S2_2/carry [19]), .B(n66508), .Q(N1319) );
  XOR21 U72946 ( .A(\sub_157_S2_2/carry [20]), .B(n66617), .Q(N1863) );
  XOR21 U72947 ( .A(\sub_126_S2_2/carry [21]), .B(n66506), .Q(N1321) );
  XOR21 U72948 ( .A(\sub_126_S2_2/carry [12]), .B(n66517), .Q(N1312) );
  XOR21 U72949 ( .A(\sub_126_S2_2/carry [14]), .B(n66515), .Q(N1314) );
  XOR21 U72950 ( .A(\sub_126_S2_2/carry [17]), .B(n66510), .Q(N1317) );
  XOR21 U72951 ( .A(\sub_126_S2_2/carry [16]), .B(n66512), .Q(N1316) );
  XOR21 U72952 ( .A(\sub_126_S2_2/carry [26]), .B(n66499), .Q(N1326) );
  XOR21 U72953 ( .A(\sub_126_S2_2/carry [28]), .B(n66497), .Q(N1328) );
  XOR21 U72954 ( .A(\sub_126_S2_2/carry [6]), .B(n66523), .Q(N1306) );
  XOR21 U72955 ( .A(\sub_157_S2_2/carry [13]), .B(n66610), .Q(N1856) );
  XOR21 U72956 ( .A(\sub_157_S2_2/carry [18]), .B(n66615), .Q(N1861) );
  XOR21 U72957 ( .A(\sub_157_S2_2/carry [27]), .B(n66625), .Q(N1870) );
  XOR21 U72958 ( .A(\sub_157_S2_2/carry [7]), .B(n66602), .Q(N1850) );
  XOR21 U72959 ( .A(\sub_126_S2_2/carry [8]), .B(n66521), .Q(N1308) );
  XOR21 U72960 ( .A(\sub_126_S2_2/carry [30]), .B(n66493), .Q(N1330) );
  XOR21 U72961 ( .A(\sub_126_S2_2/carry [4]), .B(n66525), .Q(N1304) );
  XOR21 U72962 ( .A(\sub_126_S2_2/carry [22]), .B(n66505), .Q(N1322) );
  XOR21 U72963 ( .A(\sub_157_S2_2/carry [19]), .B(n66616), .Q(N1862) );
  XOR21 U72964 ( .A(\sub_157_S2_2/carry [21]), .B(n66619), .Q(N1864) );
  XOR21 U72965 ( .A(\sub_126_S2_2/carry [15]), .B(n66514), .Q(N1315) );
  XOR21 U72966 ( .A(\sub_126_S2_2/carry [5]), .B(n66524), .Q(N1305) );
  XOR21 U72967 ( .A(\sub_126_S2_2/carry [29]), .B(n66496), .Q(N1329) );
  XOR21 U72968 ( .A(\sub_126_S2_2/carry [9]), .B(n66520), .Q(N1309) );
  XOR21 U72969 ( .A(\sub_157_S2_2/carry [12]), .B(n66609), .Q(N1855) );
  XOR21 U72970 ( .A(\sub_157_S2_2/carry [14]), .B(n66611), .Q(N1857) );
  XOR21 U72971 ( .A(\sub_157_S2_2/carry [17]), .B(n66614), .Q(N1860) );
  XOR21 U72972 ( .A(\sub_157_S2_2/carry [16]), .B(n66613), .Q(N1859) );
  XOR21 U72973 ( .A(\sub_157_S2_2/carry [26]), .B(n66624), .Q(N1869) );
  XOR21 U72974 ( .A(\sub_157_S2_2/carry [28]), .B(n66626), .Q(N1871) );
  XOR21 U72975 ( .A(\sub_157_S2_2/carry [6]), .B(n66601), .Q(N1849) );
  XOR21 U72976 ( .A(\sub_157_S2_2/carry [8]), .B(n66603), .Q(N1851) );
  XOR21 U72977 ( .A(\sub_157_S2_2/carry [30]), .B(n66583), .Q(N1873) );
  XOR21 U72978 ( .A(\sub_157_S2_2/carry [4]), .B(n66599), .Q(N1847) );
  XOR21 U72979 ( .A(\sub_157_S2_2/carry [5]), .B(n66600), .Q(N1848) );
  XOR21 U72980 ( .A(\sub_157_S2_2/carry [22]), .B(n66620), .Q(N1865) );
  XOR21 U72981 ( .A(\sub_157_S2_2/carry [15]), .B(n66612), .Q(N1858) );
  XOR21 U72982 ( .A(\sub_157_S2_2/carry [29]), .B(n66627), .Q(N1872) );
  XOR21 U72983 ( .A(\sub_157_S2_2/carry [9]), .B(n66604), .Q(N1852) );
  MUX22 U72984 ( .A(n66544), .B(n66659), .S(n65609), .Q(N3638) );
  NAND22 U72985 ( .A(n65585), .B(N3637), .Q(n66659) );
  INV3 U72986 ( .A(n66659), .Q(n66544) );
  MUX22 U72987 ( .A(n66543), .B(n66658), .S(n65609), .Q(N3511) );
  NAND22 U72988 ( .A(n65580), .B(N3510), .Q(n66658) );
  INV3 U72989 ( .A(n66658), .Q(n66543) );
  NOR31 U72990 ( .A(n66597), .B(n65545), .C(n66596), .Q(n3641) );
  XNR21 U72991 ( .A(\sub_174_2_cf/carry [4]), .B(N2052), .Q(N2072) );
  XNR21 U72992 ( .A(\sub_143_2_cf/carry[4] ), .B(N1509), .Q(N1529) );
  XNR21 U72993 ( .A(\sub_126_S2_2/carry [3]), .B(n66526), .Q(N1303) );
  XNR21 U72994 ( .A(\sub_157_S2_2/carry [3]), .B(n66598), .Q(N1846) );
  NAND22 U72995 ( .A(N2058), .B(n65740), .Q(n3375) );
  NAND22 U72996 ( .A(n3654), .B(n3364), .Q(n3425) );
  XOR21 U72997 ( .A(n65742), .B(N1506), .Q(N1526) );
  NAND22 U72998 ( .A(n3656), .B(n3358), .Q(n3415) );
  XNR21 U72999 ( .A(N4602), .B(n65580), .Q(N3359) );
  XNR21 U73000 ( .A(N4602), .B(n65585), .Q(N4605) );
  XNR21 U73001 ( .A(N4602), .B(n65583), .Q(N4468) );
  XNR21 U73002 ( .A(n65608), .B(n65578), .Q(N4329) );
  XNR21 U73003 ( .A(n65605), .B(n65578), .Q(N3377) );
  XNR21 U73004 ( .A(n65607), .B(n65578), .Q(N3204) );
  XNR21 U73005 ( .A(n65608), .B(n65578), .Q(N4730) );
  XNR21 U73006 ( .A(n65607), .B(n65578), .Q(N4456) );
  XNR21 U73007 ( .A(n65605), .B(n65578), .Q(N4593) );
  XNR21 U73008 ( .A(n66564), .B(n65582), .Q(N4190) );
  XNR21 U73009 ( .A(n66564), .B(n65585), .Q(N4317) );
  XNR21 U73010 ( .A(n66564), .B(n65583), .Q(N4857) );
  XNR21 U73011 ( .A(n66564), .B(n65580), .Q(N3395) );
  XNR21 U73012 ( .A(n66564), .B(n65584), .Q(N3222) );
  XNR21 U73013 ( .A(n66564), .B(n65585), .Q(N3049) );
  XNR21 U73014 ( .A(n66564), .B(n65583), .Q(N4718) );
  XNR21 U73015 ( .A(n66564), .B(n65583), .Q(N4581) );
  XNR21 U73016 ( .A(n66564), .B(n65584), .Q(N4444) );
  NOR31 U73017 ( .A(n66594), .B(n66597), .C(n66596), .Q(n3594) );
  NOR21 U73018 ( .A(n3601), .B(N1560), .Q(n3494) );
  XOR21 U73019 ( .A(N2049), .B(N2050), .Q(N2070) );
  NAND22 U73020 ( .A(n3711), .B(n66526), .Q(n3639) );
  NAND22 U73021 ( .A(n65740), .B(n66372), .Q(n3412) );
  NAND22 U73022 ( .A(n3586), .B(n3364), .Q(n3391) );
  XOR21 U73023 ( .A(\sub_174_2_cf/carry [3]), .B(N2051), .Q(N2071) );
  XOR21 U73024 ( .A(\sub_143_2_cf/carry[3] ), .B(N1508), .Q(N1528) );
  XOR21 U73025 ( .A(\sub_143_2_cf/carry[2] ), .B(N1507), .Q(N1527) );
  NAND22 U73026 ( .A(N1515), .B(n65741), .Q(n3350) );
  NAND22 U73027 ( .A(n3654), .B(n3489), .Q(n3419) );
  NAND22 U73028 ( .A(n65740), .B(N2049), .Q(n3397) );
  NAND22 U73029 ( .A(n65419), .B(N2049), .Q(n3411) );
  IMUX21 U73030 ( .A(n66660), .B(n66545), .S(n65609), .Q(N3900) );
  INV3 U73031 ( .A(n66660), .Q(n66545) );
  NAND22 U73032 ( .A(n65583), .B(N3899), .Q(n66660) );
  NAND22 U73033 ( .A(n3586), .B(n3489), .Q(n3438) );
  INV6 U73034 ( .A(n65595), .Q(n65594) );
  INV3 U73035 ( .A(n65596), .Q(n65593) );
  NAND22 U73036 ( .A(n3654), .B(n3473), .Q(n3511) );
  NAND22 U73037 ( .A(n3587), .B(n3494), .Q(n3389) );
  NAND22 U73038 ( .A(n3654), .B(n3456), .Q(n3506) );
  NAND22 U73039 ( .A(n65741), .B(n66539), .Q(n3407) );
  NAND22 U73040 ( .A(N1526), .B(n65742), .Q(n3372) );
  NAND22 U73041 ( .A(n65451), .B(n65740), .Q(n3352) );
  BUF6 U73042 ( .A(N690), .Q(n65936) );
  BUF6 U73043 ( .A(N684), .Q(n65946) );
  NAND41 U73044 ( .A(n66386), .B(n66331), .C(n66326), .D(n66322), .Q(n1692) );
  INV3 U73045 ( .A(n2443), .Q(n66322) );
  NAND41 U73046 ( .A(n66318), .B(n65443), .C(n66327), .D(n66390), .Q(n2244) );
  INV3 U73047 ( .A(n2273), .Q(n66390) );
  INV3 U73048 ( .A(n2315), .Q(n66327) );
  NAND41 U73049 ( .A(n66320), .B(n66329), .C(n66328), .D(n66389), .Q(n1703) );
  INV3 U73050 ( .A(n3121), .Q(n66389) );
  INV3 U73051 ( .A(n3163), .Q(n66328) );
  NAND41 U73052 ( .A(n65439), .B(n66330), .C(n66325), .D(n66321), .Q(n1730) );
  INV3 U73053 ( .A(n1931), .Q(n66321) );
  OAI2111 U73054 ( .A(n66368), .B(n66472), .C(n3603), .D(n3604), .Q(n3599) );
  INV3 U73055 ( .A(n3605), .Q(n66368) );
  NAND31 U73056 ( .A(n3594), .B(n3473), .C(n3586), .Q(n3603) );
  NAND31 U73057 ( .A(n3383), .B(n66468), .C(n3587), .Q(n3604) );
  OAI2111 U73058 ( .A(n66365), .B(n66472), .C(n3688), .D(n3689), .Q(n3680) );
  INV3 U73059 ( .A(n3706), .Q(n66365) );
  NAND31 U73060 ( .A(n3494), .B(n3561), .C(n65551), .Q(n3689) );
  NAND31 U73061 ( .A(n3364), .B(n3563), .C(n3562), .Q(n3688) );
  OAI2111 U73062 ( .A(n66367), .B(n66472), .C(n3631), .D(n3632), .Q(n3626) );
  INV3 U73063 ( .A(n3633), .Q(n66367) );
  NAND31 U73064 ( .A(n3563), .B(n3531), .C(n3364), .Q(n3631) );
  NAND31 U73065 ( .A(n3561), .B(n65548), .C(n3494), .Q(n3632) );
  OAI2111 U73066 ( .A(n66366), .B(n66472), .C(n3647), .D(n3648), .Q(n3644) );
  INV3 U73067 ( .A(n3651), .Q(n66366) );
  NAND31 U73068 ( .A(n3587), .B(n66468), .C(n65552), .Q(n3648) );
  NAND31 U73069 ( .A(n3586), .B(n3473), .C(n3641), .Q(n3647) );
  NAND41 U73070 ( .A(n66387), .B(n65439), .C(n66330), .D(n66325), .Q(n1708) );
  INV3 U73071 ( .A(n2230), .Q(n66387) );
  NAND41 U73072 ( .A(n66388), .B(n66386), .C(n66331), .D(n66326), .Q(n2413) );
  INV3 U73073 ( .A(n2780), .Q(n66388) );
  INV3 U73074 ( .A(n65611), .Q(n65610) );
  INV3 U73075 ( .A(n66871), .Q(\sub_1_root_sub_0_root_sub_167_2/A[4] ) );
  XOR21 U73076 ( .A(n65594), .B(n65585), .Q(N1120) );
  NOR21 U73077 ( .A(n66485), .B(n66395), .Q(n3380) );
  INV3 U73078 ( .A(n3587), .Q(n66485) );
  INV3 U73079 ( .A(n65920), .Q(n65915) );
  INV6 U73080 ( .A(n65920), .Q(n65918) );
  INV6 U73081 ( .A(n65580), .Q(n65578) );
  INV3 U73082 ( .A(n65546), .Q(n66537) );
  NAND31 U73083 ( .A(n3709), .B(N2046), .C(n3710), .Q(n3619) );
  NOR21 U73084 ( .A(N2063), .B(N2062), .Q(n3709) );
  NOR40 U73085 ( .A(N2067), .B(N2066), .C(N2065), .D(N2064), .Q(n3710) );
  NAND31 U73086 ( .A(n3685), .B(N1503), .C(n3686), .Q(n3615) );
  NOR21 U73087 ( .A(N1520), .B(N1519), .Q(n3685) );
  NOR40 U73088 ( .A(N1524), .B(N1523), .C(N1522), .D(N1521), .Q(n3686) );
  INV3 U73089 ( .A(n65919), .Q(n65916) );
  INV3 U73090 ( .A(n65919), .Q(n65917) );
  INV3 U73091 ( .A(n65545), .Q(n66594) );
  NOR31 U73092 ( .A(n66707), .B(n2825), .C(n66639), .Q(n2824) );
  INV3 U73093 ( .A(N3760), .Q(n66639) );
  NAND31 U73094 ( .A(N5996), .B(N5964), .C(N6028), .Q(n2825) );
  NAND31 U73095 ( .A(n66434), .B(n66383), .C(n66073), .Q(n3278) );
  INV3 U73096 ( .A(N1368), .Q(n66383) );
  INV3 U73097 ( .A(n3601), .Q(n66469) );
  NAND22 U73098 ( .A(n3656), .B(n66468), .Q(n3510) );
  INV3 U73099 ( .A(n66857), .Q(\sub_1_root_sub_0_root_sub_136_2/A[4] ) );
  NOR31 U73100 ( .A(n65425), .B(n2146), .C(n65421), .Q(n2145) );
  NAND31 U73101 ( .A(n66628), .B(N3758), .C(N3760), .Q(n2146) );
  INV3 U73102 ( .A(n3357), .Q(n66486) );
  NAND22 U73103 ( .A(n3501), .B(n66584), .Q(n3376) );
  INV3 U73104 ( .A(n3663), .Q(n66584) );
  NOR31 U73105 ( .A(n3218), .B(N1911), .C(N1914), .Q(n3279) );
  INV3 U73106 ( .A(n3344), .Q(n66472) );
  NAND22 U73107 ( .A(n3489), .B(n66576), .Q(n3333) );
  INV3 U73108 ( .A(n3381), .Q(n66535) );
  OAI2111 U73109 ( .A(n3377), .B(n66588), .C(n3433), .D(n3434), .Q(N2669) );
  AOI211 U73110 ( .A(n3437), .B(n66474), .C(n66567), .Q(n3433) );
  AOI221 U73111 ( .A(n3435), .B(n3380), .C(n65552), .D(n3382), .Q(n3434) );
  OAI2111 U73112 ( .A(n66590), .B(n3377), .C(n3378), .D(n3379), .Q(N2675) );
  AOI211 U73113 ( .A(n66474), .B(n3384), .C(n66567), .Q(n3378) );
  AOI221 U73114 ( .A(n3380), .B(n3381), .C(n3382), .D(n3383), .Q(n3379) );
  NAND22 U73115 ( .A(n3364), .B(n66576), .Q(n3342) );
  OAI2111 U73116 ( .A(n66528), .B(n3324), .C(n3325), .D(n3399), .Q(N2673) );
  AOI211 U73117 ( .A(n3337), .B(n3327), .C(n3400), .Q(n3399) );
  OAI2111 U73118 ( .A(n3324), .B(n66535), .C(n3325), .D(n3487), .Q(N2661) );
  AOI211 U73119 ( .A(n3383), .B(n3327), .C(n3488), .Q(n3487) );
  OAI2111 U73120 ( .A(n66529), .B(n3324), .C(n3325), .D(n3326), .Q(N2679) );
  AOI211 U73121 ( .A(n3327), .B(n3328), .C(n3329), .Q(n3326) );
  OAI2111 U73122 ( .A(n66529), .B(n3415), .C(n3355), .D(n3606), .Q(N2641) );
  AOI211 U73123 ( .A(n3504), .B(n3328), .C(n3607), .Q(n3606) );
  OAI2111 U73124 ( .A(n66528), .B(n3415), .C(n3355), .D(n3572), .Q(N2647) );
  AOI211 U73125 ( .A(n3504), .B(n3337), .C(n3573), .Q(n3572) );
  OAI2111 U73126 ( .A(n3415), .B(n66530), .C(n3355), .D(n3652), .Q(N2635) );
  AOI211 U73127 ( .A(n3504), .B(n3435), .C(n3653), .Q(n3652) );
  OAI2111 U73128 ( .A(n66535), .B(n66399), .C(n3325), .D(n3584), .Q(N2645) );
  AOI211 U73129 ( .A(n3380), .B(n3383), .C(n3585), .Q(n3584) );
  OAI2111 U73130 ( .A(n66535), .B(n3415), .C(n3355), .D(n3503), .Q(N2659) );
  AOI211 U73131 ( .A(n3504), .B(n3383), .C(n3505), .Q(n3503) );
  OAI2111 U73132 ( .A(n66399), .B(n66533), .C(n3325), .D(n3622), .Q(N2639) );
  AOI211 U73133 ( .A(n3562), .B(n66477), .C(n3623), .Q(n3622) );
  OAI311 U73134 ( .A(n66574), .B(n66589), .C(n66473), .D(n3624), .Q(n3623) );
  NAND31 U73135 ( .A(n3358), .B(n65548), .C(n3561), .Q(n3624) );
  OAI2111 U73136 ( .A(n66532), .B(n66399), .C(n3325), .D(n3673), .Q(N2633) );
  AOI211 U73137 ( .A(n66477), .B(n3531), .C(n3674), .Q(n3673) );
  OAI311 U73138 ( .A(n66592), .B(n66473), .C(n66574), .D(n3675), .Q(n3674) );
  NAND31 U73139 ( .A(n3561), .B(n3358), .C(n65551), .Q(n3675) );
  INV3 U73140 ( .A(n3328), .Q(n66528) );
  NAND22 U73141 ( .A(n65574), .B(n3323), .Q(n3218) );
  OAI2111 U73142 ( .A(n66589), .B(n3331), .C(n3559), .D(n3560), .Q(N2649) );
  AOI221 U73143 ( .A(n3529), .B(n65551), .C(n66397), .D(n65548), .Q(n3560) );
  AOI211 U73144 ( .A(n3530), .B(n3562), .C(n66567), .Q(n3559) );
  OAI2111 U73145 ( .A(n3331), .B(n66592), .C(n3527), .D(n3528), .Q(N2655) );
  AOI221 U73146 ( .A(n3529), .B(n65548), .C(n65551), .D(n66397), .Q(n3528) );
  AOI211 U73147 ( .A(n3530), .B(n3531), .C(n66567), .Q(n3527) );
  OAI2111 U73148 ( .A(n66473), .B(n66575), .C(n3355), .D(n3356), .Q(N2677) );
  INV3 U73149 ( .A(n3362), .Q(n66575) );
  AOI211 U73150 ( .A(n3357), .B(n3358), .C(n3359), .Q(n3356) );
  OAI2111 U73151 ( .A(n66399), .B(n66534), .C(n3325), .D(n3551), .Q(N2651) );
  AOI211 U73152 ( .A(n65552), .B(n3380), .C(n3552), .Q(n3551) );
  OAI2111 U73153 ( .A(n3415), .B(n66534), .C(n3355), .D(n3543), .Q(N2653) );
  AOI211 U73154 ( .A(n3504), .B(n65552), .C(n3544), .Q(n3543) );
  OAI2111 U73155 ( .A(n3324), .B(n66534), .C(n3325), .D(n3445), .Q(N2667) );
  AOI211 U73156 ( .A(n65552), .B(n3327), .C(n3446), .Q(n3445) );
  OAI2111 U73157 ( .A(n66533), .B(n3415), .C(n3355), .D(n3453), .Q(N2665) );
  AOI211 U73158 ( .A(n66396), .B(n65548), .C(n3454), .Q(n3453) );
  OAI2111 U73159 ( .A(n66532), .B(n3415), .C(n3355), .D(n3416), .Q(N2671) );
  AOI211 U73160 ( .A(n65551), .B(n66396), .C(n3418), .Q(n3416) );
  INV3 U73161 ( .A(n3337), .Q(n66529) );
  INV3 U73162 ( .A(n65607), .Q(n65604) );
  INV3 U73163 ( .A(n3435), .Q(n66534) );
  INV3 U73164 ( .A(n3274), .Q(n66568) );
  NOR21 U73165 ( .A(n65590), .B(n66467), .Q(n3287) );
  NAND22 U73166 ( .A(n66872), .B(n66646), .Q(n66873) );
  NAND22 U73167 ( .A(n66858), .B(n66481), .Q(n66859) );
  NOR21 U73168 ( .A(n66395), .B(n3490), .Q(n3327) );
  NAND22 U73169 ( .A(n3494), .B(n66491), .Q(n3340) );
  INV3 U73170 ( .A(n3490), .Q(n66491) );
  NAND22 U73171 ( .A(n3455), .B(n3456), .Q(n3361) );
  NAND22 U73172 ( .A(n3455), .B(n3473), .Q(n3368) );
  INV3 U73173 ( .A(N2848), .Q(n66393) );
  INV3 U73174 ( .A(n1683), .Q(n66394) );
  NAND22 U73175 ( .A(n3687), .B(n66598), .Q(n3640) );
  INV3 U73176 ( .A(n3384), .Q(n66587) );
  NAND22 U73177 ( .A(n3707), .B(\sub_174_2_cf/carry [6]), .Q(n3621) );
  NOR31 U73178 ( .A(N2046), .B(n65446), .C(N2073), .Q(n3707) );
  XNR21 U73179 ( .A(\sub_174_2_cf/carry [5]), .B(N2053), .Q(N2073) );
  NAND22 U73180 ( .A(n3683), .B(\sub_143_2_cf/carry[6] ), .Q(n3617) );
  NOR31 U73181 ( .A(N1503), .B(n65448), .C(N1530), .Q(n3683) );
  XNR21 U73182 ( .A(\sub_143_2_cf/carry[5] ), .B(N1510), .Q(N1530) );
  INV3 U73183 ( .A(N2718), .Q(n66381) );
  OAI311 U73184 ( .A(n66871), .B(n65522), .C(n3271), .D(n3275), .Q(N2718) );
  AOI311 U73185 ( .A(n3273), .B(n65742), .C(
        \sub_1_root_sub_0_root_sub_136_2/A[4] ), .D(n65547), .Q(n3275) );
  INV3 U73186 ( .A(N2719), .Q(n66382) );
  OAI311 U73187 ( .A(n66871), .B(n3271), .C(n65740), .D(n3272), .Q(N2719) );
  AOI311 U73188 ( .A(n65532), .B(n3273), .C(
        \sub_1_root_sub_0_root_sub_136_2/A[4] ), .D(n65547), .Q(n3272) );
  INV3 U73189 ( .A(n3437), .Q(n66591) );
  NAND22 U73190 ( .A(n65583), .B(N4329), .Q(n66667) );
  NAND22 U73191 ( .A(n65584), .B(N3377), .Q(n66656) );
  NAND22 U73192 ( .A(n65580), .B(N3204), .Q(n66653) );
  NAND22 U73193 ( .A(n65580), .B(N4730), .Q(n66675) );
  NAND22 U73194 ( .A(n65583), .B(N4456), .Q(n66669) );
  NAND22 U73195 ( .A(n65582), .B(N4593), .Q(n66672) );
  NAND31 U73196 ( .A(n66385), .B(n1696), .C(n66324), .Q(n1693) );
  NAND31 U73197 ( .A(n65441), .B(n1696), .C(n66323), .Q(n1731) );
  NOR21 U73198 ( .A(n2911), .B(n66697), .Q(n2910) );
  NAND31 U73199 ( .A(N5869), .B(N5837), .C(N5901), .Q(n2911) );
  NAND31 U73200 ( .A(n66323), .B(n65441), .C(n66332), .Q(n1709) );
  INV3 U73201 ( .A(n1803), .Q(n66332) );
  NAND31 U73202 ( .A(n66324), .B(n66385), .C(n66333), .Q(n2414) );
  INV3 U73203 ( .A(n2528), .Q(n66333) );
  NAND22 U73204 ( .A(n66489), .B(n66468), .Q(n3367) );
  INV3 U73205 ( .A(N2714), .Q(n66377) );
  OAI311 U73206 ( .A(n3280), .B(n65510), .C(n66871), .D(n3283), .Q(N2714) );
  AOI311 U73207 ( .A(\sub_1_root_sub_0_root_sub_136_2/A[4] ), .B(n65741), .C(
        n3282), .D(n65547), .Q(n3283) );
  INV3 U73208 ( .A(N2715), .Q(n66378) );
  OAI311 U73209 ( .A(n3280), .B(n65740), .C(n66871), .D(n3281), .Q(N2715) );
  AOI311 U73210 ( .A(\sub_1_root_sub_0_root_sub_136_2/A[4] ), .B(n65533), .C(
        n3282), .D(n65547), .Q(n3281) );
  INV3 U73211 ( .A(N2716), .Q(n66379) );
  OAI311 U73212 ( .A(n3271), .B(\sub_1_root_sub_0_root_sub_167_2/A[4] ), .C(
        n65522), .D(n3277), .Q(N2716) );
  AOI311 U73213 ( .A(n65741), .B(n66857), .C(n3273), .D(n65547), .Q(n3277) );
  INV3 U73214 ( .A(N2713), .Q(n66376) );
  OAI311 U73215 ( .A(n3280), .B(\sub_1_root_sub_0_root_sub_167_2/A[4] ), .C(
        n65740), .D(n3284), .Q(N2713) );
  AOI311 U73216 ( .A(n65533), .B(n66857), .C(n3282), .D(n65547), .Q(n3284) );
  INV3 U73217 ( .A(N2680), .Q(n66375) );
  OAI311 U73218 ( .A(n3280), .B(\sub_1_root_sub_0_root_sub_167_2/A[4] ), .C(
        n65520), .D(n3319), .Q(N2680) );
  AOI311 U73219 ( .A(n65741), .B(n66857), .C(n3282), .D(n65547), .Q(n3319) );
  NOR21 U73220 ( .A(n66490), .B(n3668), .Q(n3461) );
  INV3 U73221 ( .A(n3495), .Q(n66490) );
  INV3 U73222 ( .A(n3562), .Q(n66592) );
  INV3 U73223 ( .A(N2717), .Q(n66380) );
  OAI311 U73224 ( .A(n65740), .B(\sub_1_root_sub_0_root_sub_167_2/A[4] ), .C(
        n3271), .D(n3276), .Q(N2717) );
  AOI311 U73225 ( .A(n3273), .B(n66857), .C(n65532), .D(n65547), .Q(n3276) );
  INV3 U73226 ( .A(n3531), .Q(n66589) );
  INV3 U73227 ( .A(n66066), .Q(N1378) );
  INV3 U73228 ( .A(n66068), .Q(N1380) );
  INV3 U73229 ( .A(n66076), .Q(N1921) );
  INV3 U73230 ( .A(n66078), .Q(N1923) );
  AOI221 U73231 ( .A(n3344), .B(n3498), .C(n66469), .D(n3499), .Q(n3497) );
  AOI221 U73232 ( .A(n3344), .B(n3451), .C(n66469), .D(n3452), .Q(n3450) );
  AOI221 U73233 ( .A(n3344), .B(n3405), .C(n66469), .D(n3406), .Q(n3404) );
  AOI221 U73234 ( .A(n3344), .B(n3345), .C(n66469), .D(n3346), .Q(n3343) );
  AOI221 U73235 ( .A(n3344), .B(n3569), .C(n66469), .D(n3570), .Q(n3568) );
  AOI221 U73236 ( .A(n3344), .B(n3537), .C(n66469), .D(n3538), .Q(n3536) );
  NOR21 U73237 ( .A(n2103), .B(n65429), .Q(n2102) );
  NAND31 U73238 ( .A(N3631), .B(N3599), .C(n66636), .Q(n2103) );
  AOI221 U73239 ( .A(n65549), .B(n3592), .C(n66469), .D(n3593), .Q(n3591) );
  AOI221 U73240 ( .A(n65549), .B(n3557), .C(n66469), .D(n3558), .Q(n3556) );
  AOI221 U73241 ( .A(n65549), .B(n3521), .C(n66469), .D(n3522), .Q(n3520) );
  AOI221 U73242 ( .A(n65549), .B(n3481), .C(n66469), .D(n3482), .Q(n3480) );
  AOI221 U73243 ( .A(n65549), .B(n3443), .C(n66469), .D(n3444), .Q(n3442) );
  AOI221 U73244 ( .A(n65549), .B(n3393), .C(n66469), .D(n3394), .Q(n3392) );
  AOI221 U73245 ( .A(n65549), .B(n3661), .C(n66469), .D(n3662), .Q(n3660) );
  AOI221 U73246 ( .A(n65550), .B(n3612), .C(n66469), .D(n3613), .Q(n3611) );
  AOI221 U73247 ( .A(n65550), .B(n3578), .C(n66469), .D(n3579), .Q(n3577) );
  AOI221 U73248 ( .A(n65550), .B(n3549), .C(n66469), .D(n3550), .Q(n3548) );
  AOI221 U73249 ( .A(n65550), .B(n3513), .C(n66469), .D(n3514), .Q(n3512) );
  AOI221 U73250 ( .A(n65550), .B(n3463), .C(n66469), .D(n3464), .Q(n3462) );
  AOI221 U73251 ( .A(n65550), .B(n3427), .C(n66469), .D(n3428), .Q(n3426) );
  AOI221 U73252 ( .A(n65550), .B(n3370), .C(n66469), .D(n3371), .Q(n3369) );
  NOR21 U73253 ( .A(n66120), .B(n65452), .Q(\sub_174_2_cf/carry [4]) );
  INV3 U73254 ( .A(\sub_174_2_cf/carry [3]), .Q(n65452) );
  NOR21 U73255 ( .A(n66106), .B(n65455), .Q(\sub_143_2_cf/carry[4] ) );
  INV3 U73256 ( .A(\sub_143_2_cf/carry[3] ), .Q(n65455) );
  NOR21 U73257 ( .A(n66119), .B(n65451), .Q(\sub_174_2_cf/carry [3]) );
  INV3 U73258 ( .A(N2049), .Q(n65451) );
  NOR21 U73259 ( .A(N1361), .B(n65483), .Q(\sub_126_S2_2/carry [3]) );
  INV3 U73260 ( .A(\sub_126_S2_2/carry [2]), .Q(n65483) );
  NOR21 U73261 ( .A(n2231), .B(n65430), .Q(n2230) );
  NAND31 U73262 ( .A(N4020), .B(N3988), .C(N4021), .Q(n2231) );
  NOR21 U73263 ( .A(n2529), .B(n1805), .Q(n2528) );
  NAND31 U73264 ( .A(N7083), .B(N7051), .C(N7115), .Q(n2529) );
  NOR21 U73265 ( .A(n1804), .B(n1805), .Q(n1803) );
  NAND31 U73266 ( .A(N4813), .B(N4781), .C(N4845), .Q(n1804) );
  NOR21 U73267 ( .A(N1904), .B(n65456), .Q(\sub_157_S2_2/carry [3]) );
  INV3 U73268 ( .A(\sub_157_S2_2/carry [2]), .Q(n65456) );
  XNR21 U73269 ( .A(n65582), .B(n65603), .Q(N4041) );
  NOR21 U73270 ( .A(n2781), .B(n66631), .Q(n2780) );
  INV3 U73271 ( .A(N4021), .Q(n66631) );
  NAND31 U73272 ( .A(N6258), .B(N6226), .C(N6290), .Q(n2781) );
  NOR21 U73273 ( .A(n66105), .B(n65454), .Q(\sub_143_2_cf/carry[3] ) );
  INV3 U73274 ( .A(\sub_143_2_cf/carry[2] ), .Q(n65454) );
  NOR21 U73275 ( .A(n66104), .B(n65453), .Q(\sub_143_2_cf/carry[2] ) );
  INV3 U73276 ( .A(n65742), .Q(n65453) );
  NAND22 U73277 ( .A(n3287), .B(n3321), .Q(n3217) );
  NOR21 U73278 ( .A(N1905), .B(N1843), .Q(\sub_157_S2_2/carry [2]) );
  NOR21 U73279 ( .A(N1362), .B(N1300), .Q(\sub_126_S2_2/carry [2]) );
  NOR21 U73280 ( .A(n2274), .B(n65431), .Q(n2273) );
  NAND31 U73281 ( .A(N3040), .B(N3008), .C(n66582), .Q(n2274) );
  NOR21 U73282 ( .A(N1902), .B(n65449), .Q(\sub_157_S2_2/carry [5]) );
  NAND22 U73283 ( .A(n66489), .B(n66398), .Q(n3360) );
  INV3 U73284 ( .A(n3323), .Q(n66572) );
  NOR21 U73285 ( .A(N1359), .B(n65450), .Q(\sub_126_S2_2/carry [5]) );
  NOR21 U73286 ( .A(N1896), .B(n65462), .Q(\sub_157_S2_2/carry [11]) );
  INV3 U73287 ( .A(\sub_157_S2_2/carry [10]), .Q(n65462) );
  NOR21 U73288 ( .A(N1353), .B(n65489), .Q(\sub_126_S2_2/carry [11]) );
  INV3 U73289 ( .A(\sub_126_S2_2/carry [10]), .Q(n65489) );
  NOR21 U73290 ( .A(N1882), .B(n65476), .Q(\sub_157_S2_2/carry [25]) );
  INV3 U73291 ( .A(\sub_157_S2_2/carry [24]), .Q(n65476) );
  NOR21 U73292 ( .A(N1339), .B(n65503), .Q(\sub_126_S2_2/carry [25]) );
  INV3 U73293 ( .A(\sub_126_S2_2/carry [24]), .Q(n65503) );
  NOR21 U73294 ( .A(N1895), .B(n65463), .Q(\sub_157_S2_2/carry [12]) );
  INV3 U73295 ( .A(\sub_157_S2_2/carry [11]), .Q(n65463) );
  NOR21 U73296 ( .A(N1352), .B(n65490), .Q(\sub_126_S2_2/carry [12]) );
  INV3 U73297 ( .A(\sub_126_S2_2/carry [11]), .Q(n65490) );
  NOR21 U73298 ( .A(N1881), .B(n65477), .Q(\sub_157_S2_2/carry [26]) );
  INV3 U73299 ( .A(\sub_157_S2_2/carry [25]), .Q(n65477) );
  NOR21 U73300 ( .A(N1338), .B(n65504), .Q(\sub_126_S2_2/carry [26]) );
  INV3 U73301 ( .A(\sub_126_S2_2/carry [25]), .Q(n65504) );
  NOR21 U73302 ( .A(N1893), .B(n65465), .Q(\sub_157_S2_2/carry [14]) );
  INV3 U73303 ( .A(\sub_157_S2_2/carry [13]), .Q(n65465) );
  NOR21 U73304 ( .A(N1350), .B(n65492), .Q(\sub_126_S2_2/carry [14]) );
  INV3 U73305 ( .A(\sub_126_S2_2/carry [13]), .Q(n65492) );
  NOR21 U73306 ( .A(N1892), .B(n65466), .Q(\sub_157_S2_2/carry [15]) );
  INV3 U73307 ( .A(\sub_157_S2_2/carry [14]), .Q(n65466) );
  NOR21 U73308 ( .A(N1349), .B(n65493), .Q(\sub_126_S2_2/carry [15]) );
  INV3 U73309 ( .A(\sub_126_S2_2/carry [14]), .Q(n65493) );
  NOR21 U73310 ( .A(N1891), .B(n65467), .Q(\sub_157_S2_2/carry [16]) );
  INV3 U73311 ( .A(\sub_157_S2_2/carry [15]), .Q(n65467) );
  NOR21 U73312 ( .A(N1348), .B(n65494), .Q(\sub_126_S2_2/carry [16]) );
  INV3 U73313 ( .A(\sub_126_S2_2/carry [15]), .Q(n65494) );
  NOR21 U73314 ( .A(N1888), .B(n65470), .Q(\sub_157_S2_2/carry [19]) );
  INV3 U73315 ( .A(\sub_157_S2_2/carry [18]), .Q(n65470) );
  NOR21 U73316 ( .A(N1345), .B(n65497), .Q(\sub_126_S2_2/carry [19]) );
  INV3 U73317 ( .A(\sub_126_S2_2/carry [18]), .Q(n65497) );
  NOR21 U73318 ( .A(N1884), .B(n65474), .Q(\sub_157_S2_2/carry [23]) );
  INV3 U73319 ( .A(\sub_157_S2_2/carry [22]), .Q(n65474) );
  NOR21 U73320 ( .A(N1341), .B(n65501), .Q(\sub_126_S2_2/carry [23]) );
  INV3 U73321 ( .A(\sub_126_S2_2/carry [22]), .Q(n65501) );
  NOR21 U73322 ( .A(N1879), .B(n65479), .Q(\sub_157_S2_2/carry [28]) );
  INV3 U73323 ( .A(\sub_157_S2_2/carry [27]), .Q(n65479) );
  NOR21 U73324 ( .A(N1336), .B(n65506), .Q(\sub_126_S2_2/carry [28]) );
  INV3 U73325 ( .A(\sub_126_S2_2/carry [27]), .Q(n65506) );
  NOR21 U73326 ( .A(N1877), .B(n65481), .Q(\sub_157_S2_2/carry [30]) );
  INV3 U73327 ( .A(\sub_157_S2_2/carry [29]), .Q(n65481) );
  NOR21 U73328 ( .A(N1334), .B(n65508), .Q(\sub_126_S2_2/carry [30]) );
  INV3 U73329 ( .A(\sub_126_S2_2/carry [29]), .Q(n65508) );
  NOR21 U73330 ( .A(N1901), .B(n65457), .Q(\sub_157_S2_2/carry [6]) );
  INV3 U73331 ( .A(\sub_157_S2_2/carry [5]), .Q(n65457) );
  NOR21 U73332 ( .A(N1358), .B(n65484), .Q(\sub_126_S2_2/carry [6]) );
  INV3 U73333 ( .A(\sub_126_S2_2/carry [5]), .Q(n65484) );
  NOR21 U73334 ( .A(N1898), .B(n65460), .Q(\sub_157_S2_2/carry [9]) );
  INV3 U73335 ( .A(\sub_157_S2_2/carry [8]), .Q(n65460) );
  NOR21 U73336 ( .A(N1355), .B(n65487), .Q(\sub_126_S2_2/carry [9]) );
  INV3 U73337 ( .A(\sub_126_S2_2/carry [8]), .Q(n65487) );
  NOR21 U73338 ( .A(N1897), .B(n65461), .Q(\sub_157_S2_2/carry [10]) );
  INV3 U73339 ( .A(\sub_157_S2_2/carry [9]), .Q(n65461) );
  NOR21 U73340 ( .A(N1354), .B(n65488), .Q(\sub_126_S2_2/carry [10]) );
  INV3 U73341 ( .A(\sub_126_S2_2/carry [9]), .Q(n65488) );
  NOR21 U73342 ( .A(N1894), .B(n65464), .Q(\sub_157_S2_2/carry [13]) );
  INV3 U73343 ( .A(\sub_157_S2_2/carry [12]), .Q(n65464) );
  NOR21 U73344 ( .A(N1351), .B(n65491), .Q(\sub_126_S2_2/carry [13]) );
  INV3 U73345 ( .A(\sub_126_S2_2/carry [12]), .Q(n65491) );
  NOR21 U73346 ( .A(N1890), .B(n65468), .Q(\sub_157_S2_2/carry [17]) );
  INV3 U73347 ( .A(\sub_157_S2_2/carry [16]), .Q(n65468) );
  NOR21 U73348 ( .A(N1347), .B(n65495), .Q(\sub_126_S2_2/carry [17]) );
  INV3 U73349 ( .A(\sub_126_S2_2/carry [16]), .Q(n65495) );
  NOR21 U73350 ( .A(N1889), .B(n65469), .Q(\sub_157_S2_2/carry [18]) );
  INV3 U73351 ( .A(\sub_157_S2_2/carry [17]), .Q(n65469) );
  NOR21 U73352 ( .A(N1346), .B(n65496), .Q(\sub_126_S2_2/carry [18]) );
  INV3 U73353 ( .A(\sub_126_S2_2/carry [17]), .Q(n65496) );
  NOR21 U73354 ( .A(N1887), .B(n65471), .Q(\sub_157_S2_2/carry [20]) );
  INV3 U73355 ( .A(\sub_157_S2_2/carry [19]), .Q(n65471) );
  NOR21 U73356 ( .A(N1344), .B(n65498), .Q(\sub_126_S2_2/carry [20]) );
  INV3 U73357 ( .A(\sub_126_S2_2/carry [19]), .Q(n65498) );
  NOR21 U73358 ( .A(N1886), .B(n65472), .Q(\sub_157_S2_2/carry [21]) );
  INV3 U73359 ( .A(\sub_157_S2_2/carry [20]), .Q(n65472) );
  NOR21 U73360 ( .A(N1343), .B(n65499), .Q(\sub_126_S2_2/carry [21]) );
  INV3 U73361 ( .A(\sub_126_S2_2/carry [20]), .Q(n65499) );
  NOR21 U73362 ( .A(N1883), .B(n65475), .Q(\sub_157_S2_2/carry [24]) );
  INV3 U73363 ( .A(\sub_157_S2_2/carry [23]), .Q(n65475) );
  NOR21 U73364 ( .A(N1340), .B(n65502), .Q(\sub_126_S2_2/carry [24]) );
  INV3 U73365 ( .A(\sub_126_S2_2/carry [23]), .Q(n65502) );
  NOR21 U73366 ( .A(N1880), .B(n65478), .Q(\sub_157_S2_2/carry [27]) );
  INV3 U73367 ( .A(\sub_157_S2_2/carry [26]), .Q(n65478) );
  NOR21 U73368 ( .A(N1337), .B(n65505), .Q(\sub_126_S2_2/carry [27]) );
  INV3 U73369 ( .A(\sub_126_S2_2/carry [26]), .Q(n65505) );
  NOR21 U73370 ( .A(N1878), .B(n65480), .Q(\sub_157_S2_2/carry [29]) );
  INV3 U73371 ( .A(\sub_157_S2_2/carry [28]), .Q(n65480) );
  NOR21 U73372 ( .A(N1335), .B(n65507), .Q(\sub_126_S2_2/carry [29]) );
  INV3 U73373 ( .A(\sub_126_S2_2/carry [28]), .Q(n65507) );
  NOR21 U73374 ( .A(N1900), .B(n65458), .Q(\sub_157_S2_2/carry [7]) );
  INV3 U73375 ( .A(\sub_157_S2_2/carry [6]), .Q(n65458) );
  NOR21 U73376 ( .A(N1357), .B(n65485), .Q(\sub_126_S2_2/carry [7]) );
  INV3 U73377 ( .A(\sub_126_S2_2/carry [6]), .Q(n65485) );
  NOR21 U73378 ( .A(N1899), .B(n65459), .Q(\sub_157_S2_2/carry [8]) );
  INV3 U73379 ( .A(\sub_157_S2_2/carry [7]), .Q(n65459) );
  NOR21 U73380 ( .A(N1356), .B(n65486), .Q(\sub_126_S2_2/carry [8]) );
  INV3 U73381 ( .A(\sub_126_S2_2/carry [7]), .Q(n65486) );
  NOR21 U73382 ( .A(N1885), .B(n65473), .Q(\sub_157_S2_2/carry [22]) );
  INV3 U73383 ( .A(\sub_157_S2_2/carry [21]), .Q(n65473) );
  NOR21 U73384 ( .A(N1342), .B(n65500), .Q(\sub_126_S2_2/carry [22]) );
  INV3 U73385 ( .A(\sub_126_S2_2/carry [21]), .Q(n65500) );
  NAND31 U73386 ( .A(n3636), .B(n3637), .C(n3638), .Q(N2637) );
  NAND31 U73387 ( .A(n3586), .B(n3456), .C(n3641), .Q(n3637) );
  AOI311 U73388 ( .A(n3587), .B(n66398), .C(n65552), .D(n66567), .Q(n3636) );
  AOI221 U73389 ( .A(n3530), .B(n3437), .C(n3529), .D(n3435), .Q(n3638) );
  NAND31 U73390 ( .A(n3595), .B(n3596), .C(n3597), .Q(N2643) );
  NAND31 U73391 ( .A(n3594), .B(n3456), .C(n3586), .Q(n3596) );
  AOI311 U73392 ( .A(n3383), .B(n66398), .C(n3587), .D(n66567), .Q(n3595) );
  AOI221 U73393 ( .A(n3530), .B(n3384), .C(n3529), .D(n3381), .Q(n3597) );
  INV3 U73394 ( .A(n3286), .Q(n65576) );
  XOR31 U73395 ( .A(n65611), .B(N11344), .C(
        \add_0_root_add_0_root_sub_397_12_cf/carry [5]), .Q(N1140) );
  XOR31 U73396 ( .A(n65611), .B(N11530), .C(
        \add_0_root_add_0_root_sub_420_9_cf/carry [5]), .Q(N1266) );
  XOR31 U73397 ( .A(N5511), .B(N5517), .C(
        \add_0_root_sub_0_root_sub_375_7/carry [5]), .Q(N1032) );
  XOR31 U73398 ( .A(N5356), .B(N5362), .C(
        \add_0_root_sub_0_root_sub_372_8/carry [5]), .Q(N1014) );
  XOR31 U73399 ( .A(n65611), .B(N5208), .C(
        \add_0_root_sub_0_root_sub_369_9/carry [5]), .Q(N996) );
  BUF2 U73400 ( .A(n3436), .Q(n65552) );
  NOR31 U73401 ( .A(n66531), .B(N1300), .C(n66536), .Q(n3436) );
  INV3 U73402 ( .A(n3656), .Q(n66487) );
  INV3 U73403 ( .A(n65548), .Q(n66532) );
  INV3 U73404 ( .A(n65551), .Q(n66533) );
  BUF2 U73405 ( .A(N684), .Q(n65947) );
  BUF2 U73406 ( .A(N690), .Q(n65937) );
  NAND22 U73407 ( .A(n65443), .B(n66318), .Q(n1718) );
  NAND22 U73408 ( .A(n66329), .B(n66320), .Q(n2794) );
  BUF2 U73409 ( .A(n65592), .Q(n65590) );
  XOR31 U73410 ( .A(N3068), .B(N3074), .C(
        \add_0_root_sub_0_root_sub_300_5/carry [5]), .Q(N720) );
  BUF2 U73411 ( .A(n65592), .Q(n65591) );
  INV3 U73412 ( .A(n3502), .Q(n66585) );
  INV3 U73413 ( .A(n3496), .Q(n66494) );
  XOR31 U73414 ( .A(N6300), .B(N11332), .C(
        \add_0_root_add_0_root_sub_397_4_cf/carry [5]), .Q(N1128) );
  XOR31 U73415 ( .A(N6437), .B(N11368), .C(
        \add_0_root_add_0_root_sub_400_4_cf/carry [5]), .Q(N1146) );
  XOR31 U73416 ( .A(N6576), .B(N11392), .C(
        \add_0_root_add_0_root_sub_403_4_cf/carry [5]), .Q(N1164) );
  XOR31 U73417 ( .A(N4167), .B(N11380), .C(
        \add_0_root_add_0_root_sub_328_4_cf/carry [5]), .Q(N858) );
  XOR31 U73418 ( .A(N4306), .B(N11404), .C(
        \add_0_root_add_0_root_sub_331_4_cf/carry [5]), .Q(N876) );
  XOR31 U73419 ( .A(N3086), .B(N3092), .C(
        \add_0_root_sub_0_root_sub_300_8/carry [5]), .Q(N726) );
  INV3 U73420 ( .A(n65445), .Q(\sub_174_2_cf/carry [5]) );
  NOR21 U73421 ( .A(N2052), .B(\sub_174_2_cf/carry [4]), .Q(n65445) );
  INV3 U73422 ( .A(n65447), .Q(\sub_143_2_cf/carry[5] ) );
  NOR21 U73423 ( .A(N1509), .B(\sub_143_2_cf/carry[4] ), .Q(n65447) );
  XOR31 U73424 ( .A(N5338), .B(N5344), .C(
        \add_0_root_sub_0_root_sub_372_5/carry [5]), .Q(N1008) );
  XOR31 U73425 ( .A(n65611), .B(N2938), .C(
        \add_0_root_sub_0_root_sub_297_9/carry [5]), .Q(N708) );
  NAND31 U73426 ( .A(N4092), .B(n65440), .C(N4124), .Q(n65439) );
  INV3 U73427 ( .A(N2052), .Q(n66121) );
  INV3 U73428 ( .A(N1509), .Q(n66107) );
  INV3 U73429 ( .A(n65446), .Q(\sub_174_2_cf/carry [6]) );
  NOR21 U73430 ( .A(N2053), .B(\sub_174_2_cf/carry [5]), .Q(n65446) );
  INV3 U73431 ( .A(n65448), .Q(\sub_143_2_cf/carry[6] ) );
  NOR21 U73432 ( .A(N1510), .B(\sub_143_2_cf/carry[5] ), .Q(n65448) );
  INV3 U73433 ( .A(n65450), .Q(\sub_126_S2_2/carry [4]) );
  NOR21 U73434 ( .A(n66526), .B(\sub_126_S2_2/carry [3]), .Q(n65450) );
  INV3 U73435 ( .A(n65449), .Q(\sub_157_S2_2/carry [4]) );
  NOR21 U73436 ( .A(n66598), .B(\sub_157_S2_2/carry [3]), .Q(n65449) );
  BUF2 U73437 ( .A(n3332), .Q(n65553) );
  BUF2 U73438 ( .A(n3330), .Q(n65554) );
  NAND31 U73439 ( .A(N5058), .B(n65442), .C(N5090), .Q(n65441) );
  INV3 U73440 ( .A(n66803), .Q(n66638) );
  INV3 U73441 ( .A(n66697), .Q(n66636) );
  INV3 U73442 ( .A(n3240), .Q(n66309) );
  NOR40 U73443 ( .A(N1978), .B(N1977), .C(N1976), .D(N1975), .Q(n3240) );
  INV3 U73444 ( .A(n3266), .Q(n66236) );
  NOR40 U73445 ( .A(N1435), .B(N1434), .C(N1433), .D(N1432), .Q(n3266) );
  NAND31 U73446 ( .A(N3285), .B(n65444), .C(N3317), .Q(n65443) );
  INV3 U73447 ( .A(N2050), .Q(n66119) );
  INV3 U73448 ( .A(N1507), .Q(n66105) );
  INV3 U73449 ( .A(N2051), .Q(n66120) );
  INV3 U73450 ( .A(N1508), .Q(n66106) );
  BUF2 U73451 ( .A(n3335), .Q(n65570) );
  INV3 U73452 ( .A(N1506), .Q(n66104) );
  INV3 U73453 ( .A(n65580), .Q(n65579) );
  INV3 U73454 ( .A(n2654), .Q(n66326) );
  NOR21 U73455 ( .A(n2655), .B(n1975), .Q(n2654) );
  NAND31 U73456 ( .A(N6670), .B(N6638), .C(N6702), .Q(n2655) );
  INV3 U73457 ( .A(n1973), .Q(n66325) );
  NOR21 U73458 ( .A(n1974), .B(n1975), .Q(n1973) );
  NAND31 U73459 ( .A(N4400), .B(N4368), .C(N4432), .Q(n1974) );
  INV3 U73460 ( .A(n66707), .Q(n66628) );
  BUF2 U73461 ( .A(N683), .Q(n65949) );
  BUF2 U73462 ( .A(N689), .Q(n65939) );
  BUF2 U73463 ( .A(N683), .Q(n65948) );
  BUF2 U73464 ( .A(N689), .Q(n65938) );
  BUF2 U73465 ( .A(N683), .Q(n65950) );
  BUF2 U73466 ( .A(N689), .Q(n65940) );
  BUF2 U73467 ( .A(n65910), .Q(n65900) );
  BUF2 U73468 ( .A(n65909), .Q(n65905) );
  BUF2 U73469 ( .A(n65910), .Q(n65902) );
  BUF2 U73470 ( .A(n65908), .Q(n65906) );
  BUF2 U73471 ( .A(n65909), .Q(n65904) );
  BUF2 U73472 ( .A(n65910), .Q(n65901) );
  BUF2 U73473 ( .A(n65910), .Q(n65899) );
  BUF2 U73474 ( .A(n65837), .Q(n65903) );
  INV3 U73475 ( .A(N1510), .Q(n66108) );
  INV3 U73476 ( .A(N2053), .Q(n66122) );
  BUF2 U73477 ( .A(n65907), .Q(n65883) );
  BUF2 U73478 ( .A(n65871), .Q(n65907) );
  BUF2 U73479 ( .A(n65780), .Q(n65774) );
  BUF2 U73480 ( .A(n65780), .Q(n65775) );
  BUF2 U73481 ( .A(n65779), .Q(n65776) );
  BUF2 U73482 ( .A(n65779), .Q(n65777) );
  BUF2 U73483 ( .A(n65779), .Q(n65778) );
  BUF2 U73484 ( .A(N689), .Q(n65941) );
  BUF2 U73485 ( .A(N683), .Q(n65951) );
  INV3 U73486 ( .A(n3181), .Q(n66400) );
  AOI221 U73487 ( .A(N1874), .B(n65566), .C(N1331), .D(n66434), .Q(n3181) );
  INV3 U73488 ( .A(N2650), .Q(n66342) );
  AOI2111 U73489 ( .A(n3435), .B(n3386), .C(n3554), .D(n3555), .Q(n3553) );
  INV3 U73490 ( .A(N2666), .Q(n66346) );
  AOI2111 U73491 ( .A(n3435), .B(n3336), .C(n3448), .D(n3449), .Q(n3447) );
  INV3 U73492 ( .A(N2652), .Q(n66343) );
  AOI2111 U73493 ( .A(n3435), .B(n3421), .C(n3546), .D(n3547), .Q(n3545) );
  INV3 U73494 ( .A(N2656), .Q(n66354) );
  AOI2111 U73495 ( .A(n3386), .B(n3328), .C(n3518), .D(n3519), .Q(n3517) );
  INV3 U73496 ( .A(N2672), .Q(n66358) );
  AOI2111 U73497 ( .A(n3336), .B(n3328), .C(n3402), .D(n3403), .Q(n3401) );
  INV3 U73498 ( .A(N2646), .Q(n66353) );
  AOI2111 U73499 ( .A(n3421), .B(n3328), .C(n3575), .D(n3576), .Q(n3574) );
  INV3 U73500 ( .A(N2662), .Q(n66357) );
  AOI2111 U73501 ( .A(n3386), .B(n3337), .C(n3478), .D(n3479), .Q(n3477) );
  INV3 U73502 ( .A(N2678), .Q(n66361) );
  AOI2111 U73503 ( .A(n3336), .B(n3337), .C(n3338), .D(n3339), .Q(n3334) );
  INV3 U73504 ( .A(N2640), .Q(n66349) );
  AOI2111 U73505 ( .A(n3421), .B(n3337), .C(n3609), .D(n3610), .Q(n3608) );
  INV3 U73506 ( .A(N2660), .Q(n66356) );
  AOI2111 U73507 ( .A(n3381), .B(n3336), .C(n3492), .D(n3493), .Q(n3491) );
  INV3 U73508 ( .A(N2636), .Q(n66337) );
  AOI2111 U73509 ( .A(n3567), .B(n3435), .C(n3644), .D(n3645), .Q(n3643) );
  INV3 U73510 ( .A(N2644), .Q(n66352) );
  AOI2111 U73511 ( .A(n3386), .B(n3381), .C(n3589), .D(n3590), .Q(n3588) );
  INV3 U73512 ( .A(N2658), .Q(n66355) );
  AOI2111 U73513 ( .A(n3421), .B(n3381), .C(n3508), .D(n3509), .Q(n3507) );
  INV3 U73514 ( .A(N2642), .Q(n66350) );
  AOI2111 U73515 ( .A(n3567), .B(n3381), .C(n3599), .D(n3600), .Q(n3598) );
  INV3 U73516 ( .A(N2632), .Q(n66334) );
  AOI2111 U73517 ( .A(n3386), .B(n65548), .C(n3680), .D(n3681), .Q(n3678) );
  INV3 U73518 ( .A(N2676), .Q(n66360) );
  AOI2111 U73519 ( .A(n3362), .B(n3364), .C(n3365), .D(n3366), .Q(n3363) );
  INV3 U73520 ( .A(N2638), .Q(n66339) );
  AOI2111 U73521 ( .A(n65551), .B(n3386), .C(n3626), .D(n3627), .Q(n3625) );
  INV3 U73522 ( .A(N2664), .Q(n66345) );
  AOI2111 U73523 ( .A(n3421), .B(n65551), .C(n3458), .D(n3459), .Q(n3457) );
  INV3 U73524 ( .A(N2670), .Q(n66348) );
  AOI2111 U73525 ( .A(n3421), .B(n65548), .C(n3423), .D(n3424), .Q(n3420) );
  INV3 U73526 ( .A(n3212), .Q(n66431) );
  AOI221 U73527 ( .A(n65545), .B(n66478), .C(n65546), .D(n65565), .Q(n3212) );
  INV3 U73528 ( .A(N2648), .Q(n66341) );
  AOI2111 U73529 ( .A(n3336), .B(n65548), .C(n3565), .D(n3566), .Q(n3564) );
  INV3 U73530 ( .A(N2654), .Q(n66344) );
  AOI2111 U73531 ( .A(n65551), .B(n3336), .C(n3533), .D(n3534), .Q(n3532) );
  NOR40 U73532 ( .A(n3163), .B(n3121), .C(n1696), .D(n1691), .Q(n1724) );
  INV3 U73533 ( .A(n3677), .Q(n66467) );
  NAND22 U73534 ( .A(n66467), .B(n1691), .Q(n1683) );
  AOI311 U73535 ( .A(n66319), .B(n1689), .C(n1690), .D(n1691), .Q(n1688) );
  INV3 U73536 ( .A(n1703), .Q(n66319) );
  NOR31 U73537 ( .A(n2910), .B(n2780), .C(n2824), .Q(n1689) );
  NOR40 U73538 ( .A(n1692), .B(n1693), .C(n2528), .D(n2486), .Q(n1690) );
  XOR31 U73539 ( .A(N4330), .B(n65600), .C(\r31195/carry[5] ), .Q(N11410) );
  IMUX21 U73540 ( .A(n66667), .B(n66546), .S(N4728), .Q(N4330) );
  INV3 U73541 ( .A(n66667), .Q(n66546) );
  XOR31 U73542 ( .A(N4457), .B(n65600), .C(\r32996/carry [5]), .Q(N11428) );
  IMUX21 U73543 ( .A(n66669), .B(n66547), .S(N4728), .Q(N4457) );
  INV3 U73544 ( .A(n66669), .Q(n66547) );
  XOR31 U73545 ( .A(N7152), .B(n65600), .C(\add_417_5/carry[5] ), .Q(N11506)
         );
  XOR21 U73546 ( .A(n65610), .B(n66677), .Q(N7152) );
  NAND22 U73547 ( .A(n65577), .B(n65602), .Q(n66677) );
  XOR31 U73548 ( .A(N7278), .B(n65600), .C(\add_420_3/carry[5] ), .Q(N11524)
         );
  XOR21 U73549 ( .A(n65610), .B(n66680), .Q(N7278) );
  NAND22 U73550 ( .A(n65577), .B(m[1]), .Q(n66680) );
  XOR31 U73551 ( .A(N4882), .B(n65600), .C(\add_345_5/carry[5] ), .Q(N11518)
         );
  XOR21 U73552 ( .A(n65610), .B(n66676), .Q(N4882) );
  NAND22 U73553 ( .A(n65577), .B(n65604), .Q(n66676) );
  XOR31 U73554 ( .A(N5008), .B(n[5]), .C(\add_348_3/carry[5] ), .Q(N11536) );
  XOR21 U73555 ( .A(n65610), .B(n66679), .Q(N5008) );
  NAND22 U73556 ( .A(n65577), .B(m[1]), .Q(n66679) );
  NOR32 U73557 ( .A(N1362), .B(N1300), .C(n66531), .Q(n3328) );
  NAND22 U73558 ( .A(n65945), .B(n65521), .Q(n3177) );
  NAND22 U73559 ( .A(n65955), .B(n65533), .Q(n3178) );
  NOR32 U73560 ( .A(n66531), .B(N1362), .C(n66537), .Q(n3337) );
  NOR32 U73561 ( .A(n66537), .B(N1361), .C(n66536), .Q(n3435) );
  AOI211 U73562 ( .A(n65741), .B(N1293), .C(n66858), .Q(n66857) );
  NOR40 U73563 ( .A(n3012), .B(n3013), .C(n3014), .D(n3015), .Q(n3011) );
  NOR40 U73564 ( .A(n3052), .B(n3053), .C(n3054), .D(n3055), .Q(n3009) );
  NOR40 U73565 ( .A(n3032), .B(n3033), .C(n3034), .D(n3035), .Q(n3010) );
  NAND41 U73566 ( .A(n3698), .B(n3699), .C(n3700), .D(n3701), .Q(n3650) );
  NOR31 U73567 ( .A(N1889), .B(N1893), .C(N1891), .Q(n3700) );
  NOR31 U73568 ( .A(N1875), .B(N1879), .C(N1877), .Q(n3698) );
  NOR40 U73569 ( .A(N1901), .B(N1899), .C(N1897), .D(N1895), .Q(n3701) );
  NAND41 U73570 ( .A(n3712), .B(n3713), .C(n3714), .D(n3715), .Q(n3649) );
  NOR31 U73571 ( .A(N1346), .B(N1350), .C(N1348), .Q(n3714) );
  NOR31 U73572 ( .A(N1332), .B(N1336), .C(N1334), .Q(n3712) );
  NOR40 U73573 ( .A(N1358), .B(N1356), .C(N1354), .D(N1352), .Q(n3715) );
  XOR21 U73574 ( .A(\r2195/n3 ), .B(N1838), .Q(N2052) );
  XOR21 U73575 ( .A(\r2182/n3 ), .B(N1295), .Q(N1509) );
  NAND22 U73576 ( .A(n3677), .B(n3321), .Q(n3601) );
  XOR21 U73577 ( .A(n66483), .B(\sub_126_S2_2/carry [31]), .Q(N1331) );
  INV3 U73578 ( .A(N1332), .Q(n66483) );
  NOR21 U73579 ( .A(N1333), .B(n65509), .Q(\sub_126_S2_2/carry [31]) );
  INV3 U73580 ( .A(\sub_126_S2_2/carry [30]), .Q(n65509) );
  XOR21 U73581 ( .A(n66571), .B(\sub_157_S2_2/carry [31]), .Q(N1874) );
  INV3 U73582 ( .A(N1875), .Q(n66571) );
  NOR21 U73583 ( .A(N1876), .B(n65482), .Q(\sub_157_S2_2/carry [31]) );
  INV3 U73584 ( .A(\sub_157_S2_2/carry [30]), .Q(n65482) );
  INV3 U73585 ( .A(n66681), .Q(n66540) );
  NOR21 U73586 ( .A(n65741), .B(N1293), .Q(n66681) );
  INV3 U73587 ( .A(n66682), .Q(n66647) );
  NOR21 U73588 ( .A(n65740), .B(N1836), .Q(n66682) );
  XNR21 U73589 ( .A(N1836), .B(n65740), .Q(N689) );
  XNR21 U73590 ( .A(N1293), .B(n65741), .Q(N683) );
  NAND41 U73591 ( .A(N4436), .B(n66632), .C(N4434), .D(n66579), .Q(n1975) );
  INV3 U73592 ( .A(n66771), .Q(n66632) );
  NAND41 U73593 ( .A(N4849), .B(n66630), .C(N4847), .D(n66579), .Q(n1805) );
  INV3 U73594 ( .A(n66813), .Q(n66630) );
  NOR40 U73595 ( .A(n66590), .B(n3376), .C(N1902), .D(N1903), .Q(n3362) );
  NAND41 U73596 ( .A(n66850), .B(n66849), .C(n66848), .D(n66847), .Q(n66856)
         );
  NAND41 U73597 ( .A(n66854), .B(n66853), .C(n66852), .D(n66851), .Q(n66855)
         );
  NOR31 U73598 ( .A(n[23]), .B(n[25]), .C(n[24]), .Q(n66850) );
  NAND41 U73599 ( .A(n66721), .B(n66720), .C(n66719), .D(n66718), .Q(n66727)
         );
  NAND41 U73600 ( .A(n66725), .B(n66724), .C(n66723), .D(n66722), .Q(n66726)
         );
  NOR31 U73601 ( .A(n[23]), .B(n[25]), .C(n[24]), .Q(n66721) );
  NAND41 U73602 ( .A(n66786), .B(n66785), .C(n66784), .D(n66783), .Q(n66792)
         );
  NAND41 U73603 ( .A(n66790), .B(n66789), .C(n66788), .D(n66787), .Q(n66791)
         );
  NOR31 U73604 ( .A(n[23]), .B(n[25]), .C(n[24]), .Q(n66786) );
  NAND41 U73605 ( .A(n66711), .B(n66710), .C(n66709), .D(n66708), .Q(n66717)
         );
  NAND41 U73606 ( .A(n66715), .B(n66714), .C(n66713), .D(n66712), .Q(n66716)
         );
  NOR31 U73607 ( .A(n65593), .B(n65600), .C(n65599), .Q(n66709) );
  NOR40 U73608 ( .A(n66527), .B(n66488), .C(N1359), .D(N1360), .Q(n3357) );
  INV3 U73609 ( .A(N1905), .Q(n66596) );
  NOR31 U73610 ( .A(n66594), .B(N1904), .C(n66596), .Q(n3437) );
  NOR31 U73611 ( .A(N1904), .B(n65545), .C(n66596), .Q(n3384) );
  AOI211 U73612 ( .A(n66706), .B(n66643), .C(n66705), .Q(n66707) );
  AOI311 U73613 ( .A(n66704), .B(n66703), .C(n66702), .D(n[31]), .Q(n66705) );
  NAND41 U73614 ( .A(n66701), .B(n66700), .C(n66699), .D(n66698), .Q(n66706)
         );
  NOR40 U73615 ( .A(n66640), .B(n[16]), .C(n[18]), .D(n[17]), .Q(n66702) );
  AOI211 U73616 ( .A(n66737), .B(n66643), .C(n66736), .Q(n66738) );
  AOI311 U73617 ( .A(n66735), .B(n66734), .C(n66733), .D(n[31]), .Q(n66736) );
  NAND41 U73618 ( .A(n66732), .B(n66731), .C(n66730), .D(n66729), .Q(n66737)
         );
  NOR31 U73619 ( .A(n[24]), .B(n[26]), .C(n[25]), .Q(n66735) );
  AOI211 U73620 ( .A(n66802), .B(n66643), .C(n66801), .Q(n66803) );
  AOI311 U73621 ( .A(n66800), .B(n66799), .C(n66798), .D(n[31]), .Q(n66801) );
  NAND41 U73622 ( .A(n66796), .B(n66795), .C(n66794), .D(n66793), .Q(n66802)
         );
  NOR31 U73623 ( .A(n[24]), .B(n[26]), .C(n[25]), .Q(n66800) );
  AOI211 U73624 ( .A(n66696), .B(n66643), .C(n66695), .Q(n66697) );
  AOI311 U73625 ( .A(n66694), .B(n66693), .C(n66692), .D(n[31]), .Q(n66695) );
  NAND41 U73626 ( .A(n66691), .B(n66690), .C(n66689), .D(n66688), .Q(n66696)
         );
  NOR31 U73627 ( .A(n[24]), .B(n[26]), .C(n[25]), .Q(n66694) );
  NOR31 U73628 ( .A(n66598), .B(N1902), .C(n3376), .Q(n3654) );
  IMUX40 U73629 ( .A(n65729), .B(\GFill[4][0] ), .C(\GFill[7][0] ), .D(
        \GFill[6][0] ), .S0(n65904), .S1(N722), .Q(n7197) );
  NOR21 U73630 ( .A(N1838), .B(n66873), .Q(N1914) );
  NOR21 U73631 ( .A(N1295), .B(n66859), .Q(N1371) );
  NOR40 U73632 ( .A(n3072), .B(n3073), .C(n3074), .D(n3075), .Q(n3008) );
  NAND31 U73633 ( .A(n3076), .B(n3077), .C(n3078), .Q(n3075) );
  NAND41 U73634 ( .A(n3089), .B(n3090), .C(n3091), .D(n3092), .Q(n3072) );
  NAND41 U73635 ( .A(n3085), .B(n3086), .C(n3087), .D(n3088), .Q(n3073) );
  INV3 U73636 ( .A(N1361), .Q(n66531) );
  NOR40 U73637 ( .A(n[13]), .B(n[12]), .C(n[11]), .D(n[10]), .Q(n66732) );
  NOR40 U73638 ( .A(n[13]), .B(n[12]), .C(n[11]), .D(n[10]), .Q(n66764) );
  NOR40 U73639 ( .A(n[13]), .B(n[12]), .C(n[11]), .D(n[10]), .Q(n66829) );
  NOR40 U73640 ( .A(n[13]), .B(n[12]), .C(n[11]), .D(n[10]), .Q(n66796) );
  NOR40 U73641 ( .A(n[13]), .B(n[12]), .C(n[11]), .D(n[10]), .Q(n66691) );
  NOR31 U73642 ( .A(n66526), .B(N1359), .C(n66488), .Q(n3656) );
  NOR21 U73643 ( .A(N1836), .B(n65740), .Q(n66872) );
  NOR21 U73644 ( .A(N1293), .B(n65741), .Q(n66858) );
  INV3 U73645 ( .A(N1362), .Q(n66536) );
  INV3 U73646 ( .A(N1360), .Q(n66526) );
  NAND41 U73647 ( .A(N1339), .B(N1337), .C(N1335), .D(N1333), .Q(n3692) );
  NAND41 U73648 ( .A(N1882), .B(N1880), .C(N1878), .D(N1876), .Q(n3696) );
  NAND41 U73649 ( .A(N1338), .B(N1336), .C(N1334), .D(N1332), .Q(n3671) );
  NAND41 U73650 ( .A(N1881), .B(N1879), .C(N1877), .D(N1875), .Q(n3666) );
  NOR40 U73651 ( .A(N1887), .B(N1885), .C(N1883), .D(N1881), .Q(n3699) );
  NOR40 U73652 ( .A(N1344), .B(N1342), .C(N1340), .D(N1338), .Q(n3713) );
  XNR21 U73653 ( .A(n66873), .B(N1838), .Q(N1911) );
  NOR40 U73654 ( .A(n[5]), .B(n65598), .C(n65593), .D(n65915), .Q(n66730) );
  NOR40 U73655 ( .A(n65601), .B(n65598), .C(n65593), .D(n65915), .Q(n66742) );
  NOR40 U73656 ( .A(n65601), .B(n65598), .C(n65593), .D(n65915), .Q(n66762) );
  NOR40 U73657 ( .A(n65601), .B(n65598), .C(n65594), .D(n65915), .Q(n66827) );
  NOR40 U73658 ( .A(n65601), .B(n65598), .C(n65594), .D(n[30]), .Q(n66837) );
  NOR40 U73659 ( .A(n65601), .B(n65598), .C(n65594), .D(n[30]), .Q(n66848) );
  NOR40 U73660 ( .A(n65601), .B(n65598), .C(n65594), .D(n65915), .Q(n66805) );
  NOR40 U73661 ( .A(n65601), .B(n65598), .C(n65593), .D(n65915), .Q(n66794) );
  NOR40 U73662 ( .A(n65601), .B(n65598), .C(n65593), .D(n65915), .Q(n66699) );
  NOR40 U73663 ( .A(n65601), .B(n65598), .C(n65594), .D(n65915), .Q(n66689) );
  NOR40 U73664 ( .A(n65601), .B(n65598), .C(n65594), .D(n[30]), .Q(n66784) );
  NOR40 U73665 ( .A(n65600), .B(n65597), .C(n65593), .D(n[30]), .Q(n66773) );
  NOR40 U73666 ( .A(n65600), .B(n65599), .C(n65593), .D(n[30]), .Q(n66719) );
  NOR40 U73667 ( .A(n[26]), .B(n[25]), .C(n[24]), .D(n[23]), .Q(n66747) );
  NOR40 U73668 ( .A(n[26]), .B(n[25]), .C(n[24]), .D(n[23]), .Q(n66810) );
  NOR40 U73669 ( .A(n[26]), .B(n[25]), .C(n[24]), .D(n[23]), .Q(n66704) );
  NOR40 U73670 ( .A(N1208), .B(n[16]), .C(n[15]), .D(n[14]), .Q(n66763) );
  NOR40 U73671 ( .A(n65757), .B(n[16]), .C(n[15]), .D(n[14]), .Q(n66828) );
  INV3 U73672 ( .A(N1903), .Q(n66598) );
  NOR40 U73673 ( .A(n[17]), .B(n[16]), .C(n[15]), .D(n[14]), .Q(n66731) );
  NOR40 U73674 ( .A(n[16]), .B(n[15]), .C(n[14]), .D(n[13]), .Q(n66757) );
  NOR40 U73675 ( .A(n[17]), .B(n[16]), .C(n[15]), .D(n[14]), .Q(n66795) );
  NOR40 U73676 ( .A(n[17]), .B(n[16]), .C(n[15]), .D(n[14]), .Q(n66690) );
  NOR40 U73677 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66743) );
  NOR40 U73678 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66753) );
  NOR40 U73679 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66778) );
  NOR40 U73680 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66841) );
  NOR40 U73681 ( .A(n[29]), .B(n[28]), .C(n[27]), .D(n[26]), .Q(n66838) );
  NOR40 U73682 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66853) );
  NOR40 U73683 ( .A(n[29]), .B(n[28]), .C(n[27]), .D(n[26]), .Q(n66849) );
  NOR40 U73684 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66806) );
  NOR40 U73685 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66700) );
  NOR40 U73686 ( .A(n[16]), .B(n[15]), .C(n[14]), .D(n[13]), .Q(n66820) );
  NOR40 U73687 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66816) );
  NOR40 U73688 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66724) );
  NOR40 U73689 ( .A(n[29]), .B(n[28]), .C(n[27]), .D(n[26]), .Q(n66720) );
  NOR40 U73690 ( .A(n[15]), .B(n[14]), .C(n[13]), .D(n[12]), .Q(n66789) );
  NOR40 U73691 ( .A(n[29]), .B(n[28]), .C(n[27]), .D(n[26]), .Q(n66785) );
  NOR40 U73692 ( .A(n[16]), .B(n[15]), .C(n[14]), .D(n[13]), .Q(n66714) );
  NOR40 U73693 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66710) );
  INV3 U73694 ( .A(N1904), .Q(n66597) );
  NAND41 U73695 ( .A(n66821), .B(n66820), .C(n66819), .D(n66818), .Q(n66822)
         );
  NOR31 U73696 ( .A(n[17]), .B(n[19]), .C(n[18]), .Q(n66819) );
  NOR31 U73697 ( .A(n[10]), .B(n[12]), .C(n[11]), .Q(n66821) );
  NOR40 U73698 ( .A(n[23]), .B(n[22]), .C(n[21]), .D(n[20]), .Q(n66818) );
  NOR40 U73699 ( .A(n[23]), .B(n[22]), .C(n[21]), .D(n[20]), .Q(n66755) );
  NOR40 U73700 ( .A(n[23]), .B(n[22]), .C(n[21]), .D(n[20]), .Q(n66712) );
  NOR40 U73701 ( .A(n[22]), .B(n[21]), .C(n[20]), .D(n[19]), .Q(n66851) );
  NOR40 U73702 ( .A(n[22]), .B(n[21]), .C(n[20]), .D(n[19]), .Q(n66722) );
  NOR40 U73703 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66729) );
  NOR40 U73704 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66741) );
  NOR40 U73705 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66761) );
  NOR40 U73706 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66826) );
  NOR40 U73707 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66751) );
  NOR40 U73708 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66836) );
  NOR40 U73709 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66847) );
  NOR40 U73710 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66804) );
  NOR40 U73711 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66793) );
  NOR40 U73712 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66698) );
  NOR40 U73713 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66688) );
  NOR40 U73714 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66718) );
  NOR40 U73715 ( .A(n[22]), .B(n[21]), .C(n[20]), .D(n[19]), .Q(n66787) );
  NOR40 U73716 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66783) );
  NOR40 U73717 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66708) );
  NOR40 U73718 ( .A(n66640), .B(n[16]), .C(n[18]), .D(n[17]), .Q(n66840) );
  NAND41 U73719 ( .A(n66780), .B(n66779), .C(n66778), .D(n66777), .Q(n66781)
         );
  NOR21 U73720 ( .A(n[11]), .B(n[10]), .Q(n66780) );
  NAND31 U73721 ( .A(n65757), .B(n65834), .C(n65915), .Q(n66779) );
  NOR40 U73722 ( .A(n66640), .B(n[16]), .C(n[18]), .D(n[17]), .Q(n66777) );
  NAND41 U73723 ( .A(n66775), .B(n66774), .C(n66773), .D(n66772), .Q(n66782)
         );
  NOR31 U73724 ( .A(n[23]), .B(n[25]), .C(n[24]), .Q(n66775) );
  NOR40 U73725 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66772) );
  NOR40 U73726 ( .A(n[29]), .B(n[28]), .C(n[27]), .D(n[26]), .Q(n66774) );
  NAND41 U73727 ( .A(n66817), .B(n66816), .C(n66815), .D(n66814), .Q(n66823)
         );
  NOR31 U73728 ( .A(n65593), .B(n65600), .C(n65597), .Q(n66815) );
  NOR31 U73729 ( .A(n[24]), .B(n[26]), .C(n[25]), .Q(n66817) );
  NOR40 U73730 ( .A(n[9]), .B(n[8]), .C(n[7]), .D(n[6]), .Q(n66814) );
  XNR21 U73731 ( .A(n66859), .B(N1295), .Q(N1368) );
  NOR40 U73732 ( .A(n[23]), .B(n[22]), .C(n[21]), .D(n[20]), .Q(n66767) );
  NOR40 U73733 ( .A(n[23]), .B(n[22]), .C(n[21]), .D(n[20]), .Q(n66831) );
  NOR40 U73734 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66734) );
  NOR40 U73735 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66746) );
  NOR40 U73736 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66809) );
  NOR40 U73737 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66799) );
  NOR40 U73738 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66703) );
  NOR40 U73739 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66693) );
  NAND31 U73740 ( .A(n3716), .B(n3717), .C(n3718), .Q(n3668) );
  NOR31 U73741 ( .A(N1345), .B(N1349), .C(N1347), .Q(n3716) );
  NOR40 U73742 ( .A(N1357), .B(N1355), .C(N1353), .D(N1351), .Q(n3717) );
  NOR40 U73743 ( .A(n66502), .B(N1333), .C(N1337), .D(N1335), .Q(n3718) );
  NOR40 U73744 ( .A(n66642), .B(n[24]), .C(n[26]), .D(n[25]), .Q(n66766) );
  INV3 U73745 ( .A(n66765), .Q(n66642) );
  NOR40 U73746 ( .A(n[30]), .B(n[29]), .C(n[28]), .D(n[27]), .Q(n66765) );
  NOR40 U73747 ( .A(n66642), .B(n[24]), .C(n[26]), .D(n[25]), .Q(n66830) );
  NOR40 U73748 ( .A(n66641), .B(n[18]), .C(n[20]), .D(n[19]), .Q(n66733) );
  NOR40 U73749 ( .A(n66641), .B(n[18]), .C(n[20]), .D(n[19]), .Q(n66798) );
  INV3 U73750 ( .A(n66797), .Q(n66641) );
  NOR31 U73751 ( .A(n[21]), .B(n[23]), .C(n[22]), .Q(n66797) );
  NOR40 U73752 ( .A(n66641), .B(n[18]), .C(n[20]), .D(n[19]), .Q(n66692) );
  NAND31 U73753 ( .A(n65548), .B(n3711), .C(N1360), .Q(n3321) );
  NAND31 U73754 ( .A(n3531), .B(n3687), .C(N1903), .Q(n3323) );
  NAND31 U73755 ( .A(n3702), .B(n3703), .C(n3704), .Q(n3663) );
  NOR31 U73756 ( .A(N1888), .B(N1892), .C(N1890), .Q(n3702) );
  NOR40 U73757 ( .A(N1900), .B(N1898), .C(N1896), .D(N1894), .Q(n3703) );
  NOR40 U73758 ( .A(n66618), .B(N1876), .C(N1880), .D(N1878), .Q(n3704) );
  NAND31 U73759 ( .A(n3495), .B(N1360), .C(n3496), .Q(n3490) );
  NOR21 U73760 ( .A(n65590), .B(n1691), .Q(n3286) );
  NAND31 U73761 ( .A(n66596), .B(n66594), .C(N1904), .Q(n3332) );
  NOR31 U73762 ( .A(n66581), .B(n2487), .C(n66803), .Q(n2486) );
  INV3 U73763 ( .A(N4709), .Q(n66581) );
  NAND31 U73764 ( .A(N6946), .B(N6914), .C(N6978), .Q(n2487) );
  AOI2111 U73765 ( .A(n65918), .B(N1208), .C(n[11]), .D(n[10]), .Q(n66854) );
  AOI2111 U73766 ( .A(n65918), .B(N1208), .C(n[11]), .D(n[10]), .Q(n66725) );
  AOI2111 U73767 ( .A(n65918), .B(N1208), .C(n[11]), .D(n[10]), .Q(n66790) );
  OAI2111 U73768 ( .A(n65554), .B(n3377), .C(n66476), .D(n3474), .Q(N2663) );
  INV3 U73769 ( .A(n3475), .Q(n66476) );
  AOI221 U73770 ( .A(n3380), .B(n3328), .C(n3382), .D(n3337), .Q(n3474) );
  OAI2111 U73771 ( .A(n65553), .B(n3377), .C(n66475), .D(n3515), .Q(N2657) );
  INV3 U73772 ( .A(n3516), .Q(n66475) );
  AOI221 U73773 ( .A(n3380), .B(n3337), .C(n3382), .D(n3328), .Q(n3515) );
  AOI2111 U73774 ( .A(n65757), .B(n65832), .C(n[11]), .D(n[10]), .Q(n66744) );
  AOI2111 U73775 ( .A(n65757), .B(n65833), .C(n[11]), .D(n[10]), .Q(n66807) );
  AOI2111 U73776 ( .A(n65757), .B(n65875), .C(n[11]), .D(n[10]), .Q(n66701) );
  NOR31 U73777 ( .A(n3668), .B(N1359), .C(n3649), .Q(n3711) );
  NOR21 U73778 ( .A(n66124), .B(n66123), .Q(N1510) );
  INV3 U73779 ( .A(\r2182/n3 ), .Q(n66123) );
  INV3 U73780 ( .A(N1295), .Q(n66124) );
  NOR21 U73781 ( .A(n66126), .B(n66125), .Q(N2053) );
  INV3 U73782 ( .A(\r2195/n3 ), .Q(n66125) );
  INV3 U73783 ( .A(N1838), .Q(n66126) );
  NOR31 U73784 ( .A(n65426), .B(n1762), .C(n65422), .Q(n1761) );
  NAND31 U73785 ( .A(N4709), .B(N4708), .C(n66638), .Q(n1762) );
  NOR31 U73786 ( .A(n66599), .B(N1903), .C(n3376), .Q(n3455) );
  NAND41 U73787 ( .A(n66839), .B(n66838), .C(n66837), .D(n66836), .Q(n66845)
         );
  NAND41 U73788 ( .A(n66843), .B(n66842), .C(n66841), .D(n66840), .Q(n66844)
         );
  NOR31 U73789 ( .A(n[23]), .B(n[25]), .C(n[24]), .Q(n66839) );
  NOR31 U73790 ( .A(n3663), .B(N1902), .C(n3650), .Q(n3687) );
  NAND41 U73791 ( .A(n66754), .B(n66753), .C(n66752), .D(n66751), .Q(n66760)
         );
  NAND41 U73792 ( .A(n66758), .B(n66757), .C(n66756), .D(n66755), .Q(n66759)
         );
  NOR31 U73793 ( .A(n65593), .B(n65600), .C(n65599), .Q(n66752) );
  NOR31 U73794 ( .A(n65427), .B(n1932), .C(n65423), .Q(n1931) );
  NAND31 U73795 ( .A(N4572), .B(N4571), .C(N4573), .Q(n1932) );
  NOR31 U73796 ( .A(n66581), .B(n2444), .C(n66633), .Q(n2443) );
  INV3 U73797 ( .A(N4573), .Q(n66633) );
  NAND31 U73798 ( .A(N6809), .B(N6777), .C(N6841), .Q(n2444) );
  NOR31 U73799 ( .A(n65428), .B(n2316), .C(n65424), .Q(n2315) );
  NAND31 U73800 ( .A(N3195), .B(N3194), .C(N3196), .Q(n2316) );
  NOR31 U73801 ( .A(n66550), .B(n3164), .C(n66578), .Q(n3163) );
  INV3 U73802 ( .A(N3195), .Q(n66550) );
  INV3 U73803 ( .A(N3196), .Q(n66578) );
  NAND31 U73804 ( .A(N5432), .B(N5400), .C(N5464), .Q(n3164) );
  INV3 U73805 ( .A(n[31]), .Q(n66643) );
  NAND31 U73806 ( .A(N1904), .B(n66596), .C(n65545), .Q(n3330) );
  AOI211 U73807 ( .A(n66749), .B(n66643), .C(n66748), .Q(n66750) );
  AOI311 U73808 ( .A(n66747), .B(n66746), .C(n66745), .D(n[31]), .Q(n66748) );
  NAND41 U73809 ( .A(n66744), .B(n66743), .C(n66742), .D(n66741), .Q(n66749)
         );
  NOR40 U73810 ( .A(n66640), .B(n[16]), .C(n[18]), .D(n[17]), .Q(n66745) );
  AOI211 U73811 ( .A(n66770), .B(n66643), .C(n66769), .Q(n66771) );
  AOI311 U73812 ( .A(n66768), .B(n66767), .C(n66766), .D(n[31]), .Q(n66769) );
  NAND41 U73813 ( .A(n66764), .B(n66763), .C(n66762), .D(n66761), .Q(n66770)
         );
  NOR31 U73814 ( .A(n[17]), .B(n[19]), .C(n[18]), .Q(n66768) );
  AOI211 U73815 ( .A(n66834), .B(n66643), .C(n66833), .Q(n66835) );
  AOI311 U73816 ( .A(n66832), .B(n66831), .C(n66830), .D(n[31]), .Q(n66833) );
  NAND41 U73817 ( .A(n66829), .B(n66828), .C(n66827), .D(n66826), .Q(n66834)
         );
  NOR31 U73818 ( .A(n[17]), .B(n[19]), .C(n[18]), .Q(n66832) );
  AOI211 U73819 ( .A(n66812), .B(n66643), .C(n66811), .Q(n66813) );
  AOI311 U73820 ( .A(n66810), .B(n66809), .C(n66808), .D(n[31]), .Q(n66811) );
  NAND41 U73821 ( .A(n66807), .B(n66806), .C(n66805), .D(n66804), .Q(n66812)
         );
  NOR40 U73822 ( .A(n66640), .B(n[16]), .C(n[18]), .D(n[17]), .Q(n66808) );
  INV3 U73823 ( .A(N1837), .Q(n66646) );
  INV3 U73824 ( .A(N1294), .Q(n66481) );
  INV3 U73825 ( .A(N1902), .Q(n66599) );
  NAND31 U73826 ( .A(n66579), .B(N3349), .C(N3351), .Q(n2358) );
  INV3 U73827 ( .A(n66686), .Q(n66579) );
  XOR31 U73828 ( .A(N3241), .B(N3247), .C(
        \add_0_root_sub_0_root_sub_303_7/carry [5]), .Q(N744) );
  NAND31 U73829 ( .A(n66582), .B(N5122), .C(N5124), .Q(n1890) );
  INV3 U73830 ( .A(n66846), .Q(n66582) );
  XOR31 U73831 ( .A(n65611), .B(N11542), .C(
        \add_0_root_add_0_root_sub_348_9_cf/carry [5]), .Q(N978) );
  NAND31 U73832 ( .A(n66582), .B(N4156), .C(n66637), .Q(n2060) );
  INV3 U73833 ( .A(n66738), .Q(n66637) );
  NOR21 U73834 ( .A(n3690), .B(n3691), .Q(n3496) );
  NAND41 U73835 ( .A(n66495), .B(N1345), .C(N1341), .D(N1343), .Q(n3691) );
  NAND41 U73836 ( .A(n66513), .B(N1359), .C(N1355), .D(N1357), .Q(n3690) );
  INV3 U73837 ( .A(n3692), .Q(n66495) );
  XNR21 U73838 ( .A(n65583), .B(n65602), .Q(N5355) );
  XNR21 U73839 ( .A(n65582), .B(n65602), .Q(N3085) );
  XNR21 U73840 ( .A(n65582), .B(n65602), .Q(N6311) );
  XNR21 U73841 ( .A(n65582), .B(n65603), .Q(N6448) );
  XNR21 U73842 ( .A(n65582), .B(n65602), .Q(N5183) );
  XNR21 U73843 ( .A(n65582), .B(n65603), .Q(N4178) );
  XNR21 U73844 ( .A(n65581), .B(n65604), .Q(N7277) );
  XNR21 U73845 ( .A(n65581), .B(n65603), .Q(N7151) );
  XNR21 U73846 ( .A(n65581), .B(n65603), .Q(N4881) );
  XNR21 U73847 ( .A(n65581), .B(n65603), .Q(N5007) );
  NOR21 U73848 ( .A(n3694), .B(n3695), .Q(n3502) );
  NAND41 U73849 ( .A(n66586), .B(N1888), .C(N1884), .D(N1886), .Q(n3695) );
  NAND41 U73850 ( .A(n66606), .B(N1902), .C(N1898), .D(N1900), .Q(n3694) );
  INV3 U73851 ( .A(n3696), .Q(n66586) );
  NOR21 U73852 ( .A(n3274), .B(n66565), .Q(n3335) );
  INV3 U73853 ( .A(n3679), .Q(n66565) );
  NOR21 U73854 ( .A(n3122), .B(n66683), .Q(n3121) );
  NAND31 U73855 ( .A(N5278), .B(N5246), .C(N5310), .Q(n3122) );
  INV3 U73856 ( .A(N1359), .Q(n66525) );
  NOR31 U73857 ( .A(n[24]), .B(n[26]), .C(n[25]), .Q(n66754) );
  NOR31 U73858 ( .A(n[24]), .B(n[26]), .C(n[25]), .Q(n66711) );
  NOR31 U73859 ( .A(n[10]), .B(n[12]), .C(n[11]), .Q(n66758) );
  NOR31 U73860 ( .A(n[10]), .B(n[12]), .C(n[11]), .Q(n66715) );
  NOR31 U73861 ( .A(N1362), .B(n65546), .C(N1361), .Q(n3422) );
  BUF2 U73862 ( .A(n3417), .Q(n65551) );
  NOR31 U73863 ( .A(N1361), .B(N1362), .C(n66537), .Q(n3417) );
  NOR21 U73864 ( .A(n3669), .B(n3670), .Q(n3495) );
  NAND41 U73865 ( .A(n66492), .B(N1344), .C(N1340), .D(N1342), .Q(n3670) );
  NAND41 U73866 ( .A(n66511), .B(N1358), .C(N1354), .D(N1356), .Q(n3669) );
  INV3 U73867 ( .A(n3671), .Q(n66492) );
  NOR31 U73868 ( .A(n[17]), .B(n[19]), .C(n[18]), .Q(n66713) );
  NOR31 U73869 ( .A(n[17]), .B(n[19]), .C(n[18]), .Q(n66756) );
  NOR31 U73870 ( .A(n[16]), .B(n[18]), .C(n[17]), .Q(n66852) );
  NOR31 U73871 ( .A(n[16]), .B(n[18]), .C(n[17]), .Q(n66723) );
  NOR31 U73872 ( .A(n[16]), .B(n[18]), .C(n[17]), .Q(n66788) );
  BUF2 U73873 ( .A(N1843), .Q(n65545) );
  NOR21 U73874 ( .A(n3664), .B(n3665), .Q(n3501) );
  NAND41 U73875 ( .A(n66577), .B(N1887), .C(N1883), .D(N1885), .Q(n3665) );
  NAND41 U73876 ( .A(n66608), .B(N1901), .C(N1897), .D(N1899), .Q(n3664) );
  INV3 U73877 ( .A(n3666), .Q(n66577) );
  XOR31 U73878 ( .A(N7013), .B(n65600), .C(\add_414_5/carry[5] ), .Q(N1230) );
  XOR31 U73879 ( .A(N4743), .B(n[5]), .C(\add_342_5/carry[5] ), .Q(N942) );
  BUF2 U73880 ( .A(n65584), .Q(n65582) );
  BUF2 U73881 ( .A(n65585), .Q(n65580) );
  BUF2 U73882 ( .A(n65584), .Q(n65583) );
  INV3 U73883 ( .A(n3285), .Q(n66466) );
  AOI221 U73884 ( .A(N2045), .B(n3286), .C(N1502), .D(n65572), .Q(n3285) );
  XOR21 U73885 ( .A(\add_168/carry [31]), .B(N1982), .Q(N2045) );
  XOR21 U73886 ( .A(\add_137/carry [31]), .B(N1439), .Q(N1502) );
  INV3 U73887 ( .A(n3296), .Q(n66457) );
  AOI221 U73888 ( .A(N2036), .B(n65575), .C(N1493), .D(n65571), .Q(n3296) );
  INV3 U73889 ( .A(n3297), .Q(n66456) );
  AOI221 U73890 ( .A(N2035), .B(n65575), .C(N1492), .D(n65571), .Q(n3297) );
  INV3 U73891 ( .A(n3298), .Q(n66455) );
  AOI221 U73892 ( .A(N2034), .B(n65575), .C(N1491), .D(n65571), .Q(n3298) );
  INV3 U73893 ( .A(n3299), .Q(n66454) );
  AOI221 U73894 ( .A(N2033), .B(n65575), .C(N1490), .D(n65571), .Q(n3299) );
  INV3 U73895 ( .A(n3300), .Q(n66453) );
  AOI221 U73896 ( .A(N2032), .B(n65575), .C(N1489), .D(n65571), .Q(n3300) );
  INV3 U73897 ( .A(n3301), .Q(n66452) );
  AOI221 U73898 ( .A(N2031), .B(n65575), .C(N1488), .D(n65571), .Q(n3301) );
  INV3 U73899 ( .A(n3302), .Q(n66451) );
  AOI221 U73900 ( .A(N2030), .B(n65575), .C(N1487), .D(n65571), .Q(n3302) );
  INV3 U73901 ( .A(n3303), .Q(n66450) );
  AOI221 U73902 ( .A(N2029), .B(n65575), .C(N1486), .D(n65572), .Q(n3303) );
  INV3 U73903 ( .A(n3304), .Q(n66449) );
  AOI221 U73904 ( .A(N2028), .B(n65575), .C(N1485), .D(n65572), .Q(n3304) );
  INV3 U73905 ( .A(n3305), .Q(n66448) );
  AOI221 U73906 ( .A(N2027), .B(n65575), .C(N1484), .D(n65572), .Q(n3305) );
  INV3 U73907 ( .A(n3306), .Q(n66447) );
  AOI221 U73908 ( .A(N2026), .B(n65575), .C(N1483), .D(n65572), .Q(n3306) );
  INV3 U73909 ( .A(n3307), .Q(n66446) );
  AOI221 U73910 ( .A(N2025), .B(n65575), .C(N1482), .D(n65572), .Q(n3307) );
  INV3 U73911 ( .A(n3308), .Q(n66445) );
  AOI221 U73912 ( .A(N2024), .B(n65574), .C(N1481), .D(n65572), .Q(n3308) );
  INV3 U73913 ( .A(n3309), .Q(n66444) );
  AOI221 U73914 ( .A(N2023), .B(n65574), .C(N1480), .D(n65572), .Q(n3309) );
  INV3 U73915 ( .A(n3310), .Q(n66443) );
  AOI221 U73916 ( .A(N2022), .B(n65574), .C(N1479), .D(n65572), .Q(n3310) );
  INV3 U73917 ( .A(n3311), .Q(n66442) );
  AOI221 U73918 ( .A(N2021), .B(n65574), .C(N1478), .D(n65572), .Q(n3311) );
  INV3 U73919 ( .A(n3312), .Q(n66441) );
  AOI221 U73920 ( .A(N2020), .B(n65574), .C(N1477), .D(n65572), .Q(n3312) );
  INV3 U73921 ( .A(n3313), .Q(n66440) );
  AOI221 U73922 ( .A(N2019), .B(n65574), .C(N1476), .D(n65572), .Q(n3313) );
  INV3 U73923 ( .A(n3314), .Q(n66439) );
  AOI221 U73924 ( .A(N2018), .B(n65574), .C(N1475), .D(n65572), .Q(n3314) );
  INV3 U73925 ( .A(n3315), .Q(n66438) );
  AOI221 U73926 ( .A(N2017), .B(n65574), .C(N1474), .D(n65572), .Q(n3315) );
  INV3 U73927 ( .A(n3316), .Q(n66437) );
  AOI221 U73928 ( .A(N2016), .B(n65574), .C(N1473), .D(n65572), .Q(n3316) );
  INV3 U73929 ( .A(n3317), .Q(n66436) );
  AOI221 U73930 ( .A(N2015), .B(n65574), .C(N1472), .D(n65572), .Q(n3317) );
  INV3 U73931 ( .A(n3318), .Q(n66435) );
  AOI221 U73932 ( .A(n66595), .B(n65574), .C(n66538), .D(n3287), .Q(n3318) );
  INV3 U73933 ( .A(N2013), .Q(n66595) );
  INV3 U73934 ( .A(N1470), .Q(n66538) );
  INV3 U73935 ( .A(n3289), .Q(n66464) );
  AOI221 U73936 ( .A(N2043), .B(n3286), .C(N1500), .D(n65571), .Q(n3289) );
  INV3 U73937 ( .A(n3290), .Q(n66463) );
  AOI221 U73938 ( .A(N2042), .B(n3286), .C(N1499), .D(n65571), .Q(n3290) );
  INV3 U73939 ( .A(n3291), .Q(n66462) );
  AOI221 U73940 ( .A(N2041), .B(n3286), .C(N1498), .D(n65571), .Q(n3291) );
  INV3 U73941 ( .A(n3292), .Q(n66461) );
  AOI221 U73942 ( .A(N2040), .B(n3286), .C(N1497), .D(n65571), .Q(n3292) );
  INV3 U73943 ( .A(n3293), .Q(n66460) );
  AOI221 U73944 ( .A(N2039), .B(n3286), .C(N1496), .D(n65571), .Q(n3293) );
  INV3 U73945 ( .A(n3294), .Q(n66459) );
  AOI221 U73946 ( .A(N2038), .B(n65574), .C(N1495), .D(n65571), .Q(n3294) );
  INV3 U73947 ( .A(n3295), .Q(n66458) );
  AOI221 U73948 ( .A(N2037), .B(n65575), .C(N1494), .D(n65571), .Q(n3295) );
  INV3 U73949 ( .A(n3288), .Q(n66465) );
  AOI221 U73950 ( .A(N2044), .B(n65574), .C(N1501), .D(n65571), .Q(n3288) );
  INV3 U73951 ( .A(n3476), .Q(n66567) );
  BUF2 U73952 ( .A(n65608), .Q(n65606) );
  BUF2 U73953 ( .A(n65584), .Q(n65581) );
  BUF2 U73954 ( .A(n65608), .Q(n65605) );
  BUF2 U73955 ( .A(n65608), .Q(n65607) );
  BUF2 U73956 ( .A(n65596), .Q(n65595) );
  INV3 U73957 ( .A(N1882), .Q(n66622) );
  INV3 U73958 ( .A(N1339), .Q(n66501) );
  INV3 U73959 ( .A(N1896), .Q(n66605) );
  INV3 U73960 ( .A(N1353), .Q(n66519) );
  INV3 U73961 ( .A(N1881), .Q(n66623) );
  INV3 U73962 ( .A(N1338), .Q(n66500) );
  INV3 U73963 ( .A(N1895), .Q(n66607) );
  INV3 U73964 ( .A(N1352), .Q(n66518) );
  BUF2 U73965 ( .A(N1300), .Q(n65546) );
  INV3 U73966 ( .A(N1888), .Q(n66615) );
  INV3 U73967 ( .A(N1345), .Q(n66509) );
  INV3 U73968 ( .A(N1884), .Q(n66620) );
  INV3 U73969 ( .A(N1341), .Q(n66505) );
  INV3 U73970 ( .A(N1892), .Q(n66611) );
  INV3 U73971 ( .A(N1349), .Q(n66515) );
  INV3 U73972 ( .A(N1893), .Q(n66610) );
  INV3 U73973 ( .A(N1350), .Q(n66516) );
  INV3 U73974 ( .A(N1879), .Q(n66625) );
  INV3 U73975 ( .A(N1336), .Q(n66498) );
  INV3 U73976 ( .A(N1877), .Q(n66627) );
  INV3 U73977 ( .A(N1334), .Q(n66496) );
  INV3 U73978 ( .A(N1891), .Q(n66612) );
  INV3 U73979 ( .A(N1348), .Q(n66514) );
  INV3 U73980 ( .A(N1897), .Q(n66604) );
  INV3 U73981 ( .A(N1354), .Q(n66520) );
  INV3 U73982 ( .A(N1889), .Q(n66614) );
  INV3 U73983 ( .A(N1346), .Q(n66510) );
  INV3 U73984 ( .A(N1880), .Q(n66624) );
  INV3 U73985 ( .A(N1337), .Q(n66499) );
  INV3 U73986 ( .A(N1883), .Q(n66621) );
  INV3 U73987 ( .A(N1340), .Q(n66503) );
  INV3 U73988 ( .A(N1898), .Q(n66603) );
  INV3 U73989 ( .A(N1355), .Q(n66521) );
  INV3 U73990 ( .A(N1886), .Q(n66617) );
  INV3 U73991 ( .A(N1343), .Q(n66507) );
  INV3 U73992 ( .A(N1878), .Q(n66626) );
  INV3 U73993 ( .A(N1335), .Q(n66497) );
  INV3 U73994 ( .A(N1894), .Q(n66609) );
  INV3 U73995 ( .A(N1351), .Q(n66517) );
  INV3 U73996 ( .A(N1901), .Q(n66600) );
  INV3 U73997 ( .A(N1358), .Q(n66524) );
  INV3 U73998 ( .A(N1887), .Q(n66616) );
  INV3 U73999 ( .A(N1344), .Q(n66508) );
  INV3 U74000 ( .A(N1890), .Q(n66613) );
  INV3 U74001 ( .A(N1347), .Q(n66512) );
  INV3 U74002 ( .A(N1885), .Q(n66619) );
  INV3 U74003 ( .A(N1342), .Q(n66506) );
  INV3 U74004 ( .A(N1899), .Q(n66602) );
  INV3 U74005 ( .A(N1356), .Q(n66522) );
  INV3 U74006 ( .A(N1876), .Q(n66583) );
  INV3 U74007 ( .A(N1333), .Q(n66493) );
  INV3 U74008 ( .A(N1900), .Q(n66601) );
  INV3 U74009 ( .A(N1357), .Q(n66523) );
  XOR31 U74010 ( .A(N4996), .B(n65600), .C(\add_348/carry[5] ), .Q(N966) );
  INV3 U74011 ( .A(n3500), .Q(n66576) );
  NAND31 U74012 ( .A(n3501), .B(N1903), .C(n3502), .Q(n3500) );
  NOR21 U74013 ( .A(n[11]), .B(n[10]), .Q(n66843) );
  XOR31 U74014 ( .A(N7266), .B(n65600), .C(\add_420/carry[5] ), .Q(N1254) );
  BUF2 U74015 ( .A(n3274), .Q(n65547) );
  INV3 U74016 ( .A(n2738), .Q(n66386) );
  NOR31 U74017 ( .A(n66728), .B(n2739), .C(n66738), .Q(n2738) );
  NAND31 U74018 ( .A(N6394), .B(N6362), .C(N6426), .Q(n2739) );
  INV3 U74019 ( .A(n2399), .Q(n66318) );
  NOR21 U74020 ( .A(n2400), .B(n65432), .Q(n2399) );
  NAND31 U74021 ( .A(N3504), .B(N3472), .C(N3505), .Q(n2400) );
  INV3 U74022 ( .A(n2952), .Q(n66320) );
  NOR21 U74023 ( .A(n2953), .B(n66581), .Q(n2952) );
  NAND31 U74024 ( .A(N5742), .B(N5710), .C(N5774), .Q(n2953) );
  INV3 U74025 ( .A(n2612), .Q(n66324) );
  NOR21 U74026 ( .A(n2613), .B(n1848), .Q(n2612) );
  NAND31 U74027 ( .A(N7222), .B(N7190), .C(N7254), .Q(n2613) );
  INV3 U74028 ( .A(n1846), .Q(n66323) );
  NOR21 U74029 ( .A(n1847), .B(n1848), .Q(n1846) );
  NAND31 U74030 ( .A(N4952), .B(N4920), .C(N4984), .Q(n1847) );
  INV3 U74031 ( .A(n2994), .Q(n66329) );
  NOR31 U74032 ( .A(n66686), .B(n2995), .C(n66551), .Q(n2994) );
  INV3 U74033 ( .A(N3351), .Q(n66551) );
  NAND31 U74034 ( .A(N5587), .B(N5555), .C(N5619), .Q(n2995) );
  BUF2 U74035 ( .A(n65742), .Q(n65741) );
  INV3 U74036 ( .A(n2570), .Q(n66385) );
  NOR31 U74037 ( .A(n66846), .B(n2571), .C(n66635), .Q(n2570) );
  INV3 U74038 ( .A(N5124), .Q(n66635) );
  NAND31 U74039 ( .A(N7360), .B(N7328), .C(N7392), .Q(n2571) );
  INV3 U74040 ( .A(N2631), .Q(n65592) );
  INV3 U74041 ( .A(n66776), .Q(n66640) );
  NOR40 U74042 ( .A(n[22]), .B(n[21]), .C(n[20]), .D(n[19]), .Q(n66776) );
  INV3 U74043 ( .A(n2696), .Q(n66331) );
  NOR21 U74044 ( .A(n2697), .B(n2018), .Q(n2696) );
  NAND31 U74045 ( .A(N6531), .B(N6499), .C(N6563), .Q(n2697) );
  INV3 U74046 ( .A(n2016), .Q(n66330) );
  NOR21 U74047 ( .A(n2017), .B(n2018), .Q(n2016) );
  NAND31 U74048 ( .A(N4261), .B(N4229), .C(N4293), .Q(n2017) );
  INV3 U74049 ( .A(n3460), .Q(n66489) );
  NAND31 U74050 ( .A(N1359), .B(n66526), .C(n3461), .Q(n3460) );
  INV3 U74051 ( .A(n3672), .Q(n66511) );
  NAND41 U74052 ( .A(N1352), .B(N1350), .C(N1348), .D(N1346), .Q(n3672) );
  INV3 U74053 ( .A(n3693), .Q(n66513) );
  NAND41 U74054 ( .A(N1353), .B(N1351), .C(N1349), .D(N1347), .Q(n3693) );
  INV3 U74055 ( .A(n3697), .Q(n66606) );
  NAND41 U74056 ( .A(N1896), .B(N1894), .C(N1892), .D(N1890), .Q(n3697) );
  INV3 U74057 ( .A(n3667), .Q(n66608) );
  NAND41 U74058 ( .A(N1895), .B(N1893), .C(N1891), .D(N1889), .Q(n3667) );
  INV3 U74059 ( .A(n3214), .Q(n66384) );
  AOI221 U74060 ( .A(N1838), .B(n66478), .C(N1295), .D(n65565), .Q(n3214) );
  INV3 U74061 ( .A(n3705), .Q(n66618) );
  NOR31 U74062 ( .A(N1884), .B(N1886), .C(N1882), .Q(n3705) );
  INV3 U74063 ( .A(n3719), .Q(n66502) );
  NOR31 U74064 ( .A(N1341), .B(N1343), .C(N1339), .Q(n3719) );
  INV3 U74065 ( .A(n3216), .Q(n66433) );
  AOI221 U74066 ( .A(N1293), .B(n65565), .C(N1836), .D(n66478), .Q(n3216) );
  BUF2 U74067 ( .A(n65920), .Q(n65919) );
  BUF2 U74068 ( .A(N1207), .Q(n65908) );
  BUF2 U74069 ( .A(N1207), .Q(n65909) );
  BUF2 U74070 ( .A(N1207), .Q(n65910) );
  INV3 U74071 ( .A(n3215), .Q(n66432) );
  AOI221 U74072 ( .A(N1294), .B(n65565), .C(N1837), .D(n66478), .Q(n3215) );
  BUF2 U74073 ( .A(n65781), .Q(n65780) );
  BUF2 U74074 ( .A(n65781), .Q(n65779) );
  INV3 U74075 ( .A(N2629), .Q(n66566) );
  NAND31 U74076 ( .A(n65592), .B(n65569), .C(n3476), .Q(N2629) );
  XOR31 U74077 ( .A(N6312), .B(N11338), .C(
        \add_0_root_add_0_root_sub_397_8_cf/carry [5]), .Q(N1134) );
  XOR21 U74078 ( .A(n65610), .B(n66662), .Q(N6312) );
  NAND22 U74079 ( .A(n65577), .B(n65604), .Q(n66662) );
  XOR31 U74080 ( .A(N6449), .B(N11374), .C(
        \add_0_root_add_0_root_sub_400_8_cf/carry [5]), .Q(N1152) );
  XOR21 U74081 ( .A(n65610), .B(n66664), .Q(N6449) );
  NAND22 U74082 ( .A(n65577), .B(m[1]), .Q(n66664) );
  XOR31 U74083 ( .A(N7140), .B(n[5]), .C(\add_417_3/carry[5] ), .Q(N1242) );
  XNR21 U74084 ( .A(m[2]), .B(n65603), .Q(N7140) );
  XOR31 U74085 ( .A(N5166), .B(N5172), .C(
        \add_0_root_sub_0_root_sub_369_3/carry [5]), .Q(N984) );
  XNR21 U74086 ( .A(n65609), .B(n65603), .Q(N5166) );
  XOR31 U74087 ( .A(N5184), .B(N5190), .C(
        \add_0_root_sub_0_root_sub_369_6/carry [5]), .Q(N990) );
  XOR21 U74088 ( .A(m[2]), .B(n66649), .Q(N5184) );
  NAND22 U74089 ( .A(n65578), .B(n65604), .Q(n66649) );
  XOR31 U74090 ( .A(n[5]), .B(N11350), .C(
        \add_0_root_add_0_root_sub_325_4_cf/carry [5]), .Q(N840) );
  XNR21 U74091 ( .A(n65610), .B(n65602), .Q(N4030) );
  XOR31 U74092 ( .A(n[5]), .B(N11356), .C(
        \add_0_root_add_0_root_sub_325_8_cf/carry [5]), .Q(N846) );
  XOR21 U74093 ( .A(n65609), .B(n66661), .Q(N4042) );
  IMUX21 U74094 ( .A(n66665), .B(n66556), .S(n65555), .Q(N4191) );
  INV3 U74095 ( .A(n66665), .Q(n66556) );
  NAND22 U74096 ( .A(n65577), .B(N4190), .Q(n66665) );
  XOR31 U74097 ( .A(N4179), .B(N11386), .C(
        \add_0_root_add_0_root_sub_328_8_cf/carry [5]), .Q(N864) );
  XOR21 U74098 ( .A(n65610), .B(n66663), .Q(N4179) );
  NAND22 U74099 ( .A(n65577), .B(m[1]), .Q(n66663) );
  IMUX21 U74100 ( .A(n66666), .B(n66557), .S(n65555), .Q(N4318) );
  INV3 U74101 ( .A(n66666), .Q(n66557) );
  NAND22 U74102 ( .A(n65577), .B(N4317), .Q(n66666) );
  IMUX21 U74103 ( .A(n66678), .B(n66563), .S(n65555), .Q(N4858) );
  INV3 U74104 ( .A(n66678), .Q(n66563) );
  XOR31 U74105 ( .A(N4870), .B(n[5]), .C(\add_345_3/carry[5] ), .Q(N954) );
  XNR21 U74106 ( .A(m[2]), .B(n65603), .Q(N4870) );
  IMUX21 U74107 ( .A(n66656), .B(n66542), .S(N4728), .Q(N3378) );
  INV3 U74108 ( .A(n66656), .Q(n66542) );
  IMUX21 U74109 ( .A(n66657), .B(n66555), .S(n65555), .Q(N3396) );
  INV3 U74110 ( .A(n66657), .Q(n66555) );
  IMUX21 U74111 ( .A(n66655), .B(n66554), .S(N4603), .Q(N3360) );
  INV3 U74112 ( .A(n66655), .Q(n66554) );
  IMUX21 U74113 ( .A(n66653), .B(n66541), .S(N4728), .Q(N3205) );
  INV3 U74114 ( .A(n66653), .Q(n66541) );
  IMUX21 U74115 ( .A(n66654), .B(n66553), .S(n65555), .Q(N3223) );
  INV3 U74116 ( .A(n66654), .Q(n66553) );
  IMUX21 U74117 ( .A(n66652), .B(n66552), .S(n65555), .Q(N3050) );
  INV3 U74118 ( .A(n66652), .Q(n66552) );
  XOR31 U74119 ( .A(n65600), .B(N2920), .C(
        \add_0_root_sub_0_root_sub_297_6/carry [5]), .Q(N702) );
  INV3 U74120 ( .A(n66167), .Q(n66168) );
  XOR21 U74121 ( .A(n65610), .B(n66648), .Q(N2914) );
  XOR31 U74122 ( .A(n[5]), .B(N2902), .C(
        \add_0_root_sub_0_root_sub_297_3/carry [5]), .Q(N696) );
  XNR21 U74123 ( .A(n65609), .B(n65602), .Q(N2896) );
  INV3 U74124 ( .A(n66169), .Q(n66170) );
  IMUX21 U74125 ( .A(n66674), .B(n66562), .S(n65555), .Q(N4719) );
  INV3 U74126 ( .A(n66674), .Q(n66562) );
  IMUX21 U74127 ( .A(n66675), .B(n66549), .S(N4728), .Q(N4731) );
  INV3 U74128 ( .A(n66675), .Q(n66549) );
  IMUX21 U74129 ( .A(n66673), .B(n66561), .S(N4603), .Q(N4606) );
  INV3 U74130 ( .A(n66673), .Q(n66561) );
  IMUX21 U74131 ( .A(n66671), .B(n66560), .S(n65555), .Q(N4582) );
  INV3 U74132 ( .A(n66671), .Q(n66560) );
  IMUX21 U74133 ( .A(n66672), .B(n66548), .S(N4728), .Q(N4594) );
  INV3 U74134 ( .A(n66672), .Q(n66548) );
  IMUX21 U74135 ( .A(n66670), .B(n66559), .S(N4603), .Q(N4469) );
  INV3 U74136 ( .A(n66670), .Q(n66559) );
  IMUX21 U74137 ( .A(n66668), .B(n66558), .S(n65555), .Q(N4445) );
  INV3 U74138 ( .A(n66668), .Q(n66558) );
  NAND22 U74139 ( .A(n65577), .B(N4444), .Q(n66668) );
  NAND22 U74140 ( .A(O_play[3]), .B(n1680), .Q(n1691) );
  AOI311 U74141 ( .A(n1685), .B(n1686), .C(n1687), .D(n1688), .Q(n1684) );
  NOR31 U74142 ( .A(n2145), .B(n1718), .C(n2102), .Q(n1686) );
  NOR40 U74143 ( .A(n1708), .B(n1709), .C(n1761), .D(n1931), .Q(n1687) );
  AOI311 U74144 ( .A(n1724), .B(n1725), .C(n1726), .D(n1727), .Q(n1723) );
  NOR31 U74145 ( .A(n2824), .B(n2794), .C(n2910), .Q(n1725) );
  NOR40 U74146 ( .A(n2413), .B(n2414), .C(n2486), .D(n2443), .Q(n1726) );
  NOR21 U74147 ( .A(n1680), .B(O_play[3]), .Q(n3677) );
  AOI311 U74148 ( .A(n65604), .B(n65579), .C(m[2]), .D(n66580), .Q(N3351) );
  INV3 U74149 ( .A(n66687), .Q(n66580) );
  NAND22 U74150 ( .A(state[1]), .B(n1654), .Q(n3476) );
  NAND41 U74151 ( .A(N4297), .B(n66629), .C(N4295), .D(N4294), .Q(n2018) );
  INV3 U74152 ( .A(n66750), .Q(n66629) );
  NAND22 U74153 ( .A(n66740), .B(n66739), .Q(N4294) );
  NAND41 U74154 ( .A(N4988), .B(n66634), .C(N4986), .D(N4985), .Q(n1848) );
  INV3 U74155 ( .A(n66835), .Q(n66634) );
  NAND22 U74156 ( .A(n66825), .B(n66824), .Q(N4985) );
  NOR40 U74157 ( .A(\Col_Fill[2][21] ), .B(\Col_Fill[2][20] ), .C(
        \Col_Fill[2][1] ), .D(\Col_Fill[2][19] ), .Q(n3060) );
  NOR40 U74158 ( .A(\Col_Fill[2][8] ), .B(\Col_Fill[2][7] ), .C(
        \Col_Fill[2][6] ), .D(\Col_Fill[2][5] ), .Q(n3064) );
  NOR40 U74159 ( .A(\Col_Fill[6][25] ), .B(\Col_Fill[6][24] ), .C(
        \Col_Fill[6][23] ), .D(\Col_Fill[6][22] ), .Q(n3020) );
  NOR40 U74160 ( .A(\Col_Fill[6][10] ), .B(\Col_Fill[6][0] ), .C(
        \Col_Fill[5][9] ), .D(\Col_Fill[5][8] ), .Q(n3016) );
  NOR40 U74161 ( .A(\Col_Fill[0][1] ), .B(\Col_Fill[0][19] ), .C(
        \Col_Fill[0][18] ), .D(\Col_Fill[0][17] ), .Q(n3081) );
  NOR40 U74162 ( .A(\Col_Fill[0][6] ), .B(\Col_Fill[0][5] ), .C(
        \Col_Fill[0][4] ), .D(\Col_Fill[0][31] ), .Q(n3085) );
  NOR40 U74163 ( .A(\Col_Fill[4][23] ), .B(\Col_Fill[4][22] ), .C(
        \Col_Fill[4][21] ), .D(\Col_Fill[4][20] ), .Q(n3040) );
  NOR40 U74164 ( .A(\Col_Fill[1][20] ), .B(\Col_Fill[1][1] ), .C(
        \Col_Fill[1][19] ), .D(\Col_Fill[1][18] ), .Q(n3089) );
  NOR40 U74165 ( .A(\Col_Fill[3][9] ), .B(\Col_Fill[3][8] ), .C(
        \Col_Fill[3][7] ), .D(\Col_Fill[3][6] ), .Q(n3036) );
  NOR40 U74166 ( .A(\Col_Fill[5][0] ), .B(\Col_Fill[4][9] ), .C(
        \Col_Fill[4][8] ), .D(\Col_Fill[4][7] ), .Q(n3044) );
  NOR40 U74167 ( .A(\Col_Fill[5][24] ), .B(\Col_Fill[5][23] ), .C(
        \Col_Fill[5][22] ), .D(\Col_Fill[5][21] ), .Q(n3048) );
  NOR40 U74168 ( .A(\Col_Fill[1][7] ), .B(\Col_Fill[1][6] ), .C(
        \Col_Fill[1][5] ), .D(\Col_Fill[1][4] ), .Q(n3056) );
  NOR40 U74169 ( .A(\Col_Fill[3][22] ), .B(\Col_Fill[3][21] ), .C(
        \Col_Fill[3][20] ), .D(\Col_Fill[3][1] ), .Q(n3068) );
  NOR40 U74170 ( .A(\Col_Fill[7][11] ), .B(\Col_Fill[7][10] ), .C(
        \Col_Fill[7][0] ), .D(\Col_Fill[6][9] ), .Q(n3024) );
  NOR40 U74171 ( .A(\Col_Fill[7][26] ), .B(\Col_Fill[7][25] ), .C(
        \Col_Fill[7][24] ), .D(\Col_Fill[7][23] ), .Q(n3028) );
  BUF6 U74172 ( .A(n[4]), .Q(n65597) );
  BUF6 U74173 ( .A(n[4]), .Q(n65598) );
  BUF6 U74174 ( .A(n[4]), .Q(n65599) );
  NAND41 U74175 ( .A(n3060), .B(n3061), .C(n3062), .D(n3063), .Q(n3054) );
  NOR40 U74176 ( .A(\Col_Fill[2][4] ), .B(\Col_Fill[2][31] ), .C(
        \Col_Fill[2][30] ), .D(\Col_Fill[2][2] ), .Q(n3063) );
  NOR40 U74177 ( .A(\Col_Fill[2][25] ), .B(\Col_Fill[2][24] ), .C(
        \Col_Fill[2][23] ), .D(\Col_Fill[2][22] ), .Q(n3061) );
  NOR40 U74178 ( .A(\Col_Fill[2][29] ), .B(\Col_Fill[2][28] ), .C(
        \Col_Fill[2][27] ), .D(\Col_Fill[2][26] ), .Q(n3062) );
  NAND41 U74179 ( .A(n3020), .B(n3021), .C(n3022), .D(n3023), .Q(n3014) );
  NOR40 U74180 ( .A(\Col_Fill[6][8] ), .B(\Col_Fill[6][7] ), .C(
        \Col_Fill[6][6] ), .D(\Col_Fill[6][5] ), .Q(n3023) );
  NOR40 U74181 ( .A(\Col_Fill[6][29] ), .B(\Col_Fill[6][28] ), .C(
        \Col_Fill[6][27] ), .D(\Col_Fill[6][26] ), .Q(n3021) );
  NOR40 U74182 ( .A(\Col_Fill[6][4] ), .B(\Col_Fill[6][31] ), .C(
        \Col_Fill[6][30] ), .D(\Col_Fill[6][2] ), .Q(n3022) );
  NAND41 U74183 ( .A(n3081), .B(n3082), .C(n3083), .D(n3084), .Q(n3074) );
  NOR40 U74184 ( .A(\Col_Fill[0][30] ), .B(\Col_Fill[0][2] ), .C(
        \Col_Fill[0][29] ), .D(\Col_Fill[0][28] ), .Q(n3084) );
  NOR40 U74185 ( .A(\Col_Fill[0][23] ), .B(\Col_Fill[0][22] ), .C(
        \Col_Fill[0][21] ), .D(\Col_Fill[0][20] ), .Q(n3082) );
  NOR40 U74186 ( .A(\Col_Fill[0][27] ), .B(\Col_Fill[0][26] ), .C(
        \Col_Fill[0][25] ), .D(\Col_Fill[0][24] ), .Q(n3083) );
  NAND41 U74187 ( .A(n3040), .B(n3041), .C(n3042), .D(n3043), .Q(n3034) );
  NOR40 U74188 ( .A(\Col_Fill[4][6] ), .B(\Col_Fill[4][5] ), .C(
        \Col_Fill[4][4] ), .D(\Col_Fill[4][31] ), .Q(n3043) );
  NOR40 U74189 ( .A(\Col_Fill[4][27] ), .B(\Col_Fill[4][26] ), .C(
        \Col_Fill[4][25] ), .D(\Col_Fill[4][24] ), .Q(n3041) );
  NOR40 U74190 ( .A(\Col_Fill[4][30] ), .B(\Col_Fill[4][2] ), .C(
        \Col_Fill[4][29] ), .D(\Col_Fill[4][28] ), .Q(n3042) );
  NAND41 U74191 ( .A(n3064), .B(n3065), .C(n3066), .D(n3067), .Q(n3053) );
  NOR40 U74192 ( .A(\Col_Fill[3][19] ), .B(\Col_Fill[3][18] ), .C(
        \Col_Fill[3][17] ), .D(\Col_Fill[3][16] ), .Q(n3067) );
  NOR40 U74193 ( .A(\Col_Fill[3][11] ), .B(\Col_Fill[3][10] ), .C(
        \Col_Fill[3][0] ), .D(\Col_Fill[2][9] ), .Q(n3065) );
  NOR40 U74194 ( .A(\Col_Fill[3][15] ), .B(\Col_Fill[3][14] ), .C(
        \Col_Fill[3][13] ), .D(\Col_Fill[3][12] ), .Q(n3066) );
  NAND41 U74195 ( .A(n3016), .B(n3017), .C(n3018), .D(n3019), .Q(n3015) );
  NOR40 U74196 ( .A(\Col_Fill[6][21] ), .B(\Col_Fill[6][20] ), .C(
        \Col_Fill[6][1] ), .D(\Col_Fill[6][19] ), .Q(n3019) );
  NOR40 U74197 ( .A(\Col_Fill[6][14] ), .B(\Col_Fill[6][13] ), .C(
        \Col_Fill[6][12] ), .D(\Col_Fill[6][11] ), .Q(n3017) );
  NOR40 U74198 ( .A(\Col_Fill[6][18] ), .B(\Col_Fill[6][17] ), .C(
        \Col_Fill[6][16] ), .D(\Col_Fill[6][15] ), .Q(n3018) );
  NAND41 U74199 ( .A(n3036), .B(n3037), .C(n3038), .D(n3039), .Q(n3035) );
  NOR40 U74200 ( .A(\Col_Fill[4][1] ), .B(\Col_Fill[4][19] ), .C(
        \Col_Fill[4][18] ), .D(\Col_Fill[4][17] ), .Q(n3039) );
  NOR40 U74201 ( .A(\Col_Fill[4][12] ), .B(\Col_Fill[4][11] ), .C(
        \Col_Fill[4][10] ), .D(\Col_Fill[4][0] ), .Q(n3037) );
  NOR40 U74202 ( .A(\Col_Fill[4][16] ), .B(\Col_Fill[4][15] ), .C(
        \Col_Fill[4][14] ), .D(\Col_Fill[4][13] ), .Q(n3038) );
  NAND41 U74203 ( .A(n3044), .B(n3045), .C(n3046), .D(n3047), .Q(n3033) );
  NOR40 U74204 ( .A(\Col_Fill[5][20] ), .B(\Col_Fill[5][1] ), .C(
        \Col_Fill[5][19] ), .D(\Col_Fill[5][18] ), .Q(n3047) );
  NOR40 U74205 ( .A(\Col_Fill[5][13] ), .B(\Col_Fill[5][12] ), .C(
        \Col_Fill[5][11] ), .D(\Col_Fill[5][10] ), .Q(n3045) );
  NOR40 U74206 ( .A(\Col_Fill[5][17] ), .B(\Col_Fill[5][16] ), .C(
        \Col_Fill[5][15] ), .D(\Col_Fill[5][14] ), .Q(n3046) );
  NAND41 U74207 ( .A(n3056), .B(n3057), .C(n3058), .D(n3059), .Q(n3055) );
  NOR40 U74208 ( .A(\Col_Fill[2][18] ), .B(\Col_Fill[2][17] ), .C(
        \Col_Fill[2][16] ), .D(\Col_Fill[2][15] ), .Q(n3059) );
  NOR40 U74209 ( .A(\Col_Fill[2][10] ), .B(\Col_Fill[2][0] ), .C(
        \Col_Fill[1][9] ), .D(\Col_Fill[1][8] ), .Q(n3057) );
  NOR40 U74210 ( .A(\Col_Fill[2][14] ), .B(\Col_Fill[2][13] ), .C(
        \Col_Fill[2][12] ), .D(\Col_Fill[2][11] ), .Q(n3058) );
  NAND41 U74211 ( .A(n3024), .B(n3025), .C(n3026), .D(n3027), .Q(n3013) );
  NOR40 U74212 ( .A(\Col_Fill[7][22] ), .B(\Col_Fill[7][21] ), .C(
        \Col_Fill[7][20] ), .D(\Col_Fill[7][1] ), .Q(n3027) );
  NOR40 U74213 ( .A(\Col_Fill[7][15] ), .B(\Col_Fill[7][14] ), .C(
        \Col_Fill[7][13] ), .D(\Col_Fill[7][12] ), .Q(n3025) );
  NOR40 U74214 ( .A(\Col_Fill[7][19] ), .B(\Col_Fill[7][18] ), .C(
        \Col_Fill[7][17] ), .D(\Col_Fill[7][16] ), .Q(n3026) );
  NOR40 U74215 ( .A(\Col_Fill[0][16] ), .B(\Col_Fill[0][15] ), .C(
        \Col_Fill[0][14] ), .D(\Col_Fill[0][13] ), .Q(n3077) );
  NAND41 U74216 ( .A(n3048), .B(n3049), .C(n3050), .D(n3051), .Q(n3032) );
  NOR40 U74217 ( .A(\Col_Fill[5][7] ), .B(\Col_Fill[5][6] ), .C(
        \Col_Fill[5][5] ), .D(\Col_Fill[5][4] ), .Q(n3051) );
  NOR40 U74218 ( .A(\Col_Fill[5][28] ), .B(\Col_Fill[5][27] ), .C(
        \Col_Fill[5][26] ), .D(\Col_Fill[5][25] ), .Q(n3049) );
  NOR40 U74219 ( .A(\Col_Fill[5][31] ), .B(\Col_Fill[5][30] ), .C(
        \Col_Fill[5][2] ), .D(\Col_Fill[5][29] ), .Q(n3050) );
  NAND41 U74220 ( .A(n3068), .B(n3069), .C(n3070), .D(n3071), .Q(n3052) );
  NOR40 U74221 ( .A(\Col_Fill[3][5] ), .B(\Col_Fill[3][4] ), .C(
        \Col_Fill[3][31] ), .D(\Col_Fill[3][30] ), .Q(n3071) );
  NOR40 U74222 ( .A(\Col_Fill[3][26] ), .B(\Col_Fill[3][25] ), .C(
        \Col_Fill[3][24] ), .D(\Col_Fill[3][23] ), .Q(n3069) );
  NOR40 U74223 ( .A(\Col_Fill[3][2] ), .B(\Col_Fill[3][29] ), .C(
        \Col_Fill[3][28] ), .D(\Col_Fill[3][27] ), .Q(n3070) );
  NAND41 U74224 ( .A(n3028), .B(n3029), .C(n3030), .D(n3031), .Q(n3012) );
  NOR40 U74225 ( .A(\Col_Fill[7][9] ), .B(\Col_Fill[7][8] ), .C(
        \Col_Fill[7][7] ), .D(\Col_Fill[7][6] ), .Q(n3031) );
  NOR40 U74226 ( .A(\Col_Fill[7][2] ), .B(\Col_Fill[7][29] ), .C(
        \Col_Fill[7][28] ), .D(\Col_Fill[7][27] ), .Q(n3029) );
  NOR40 U74227 ( .A(\Col_Fill[7][5] ), .B(\Col_Fill[7][4] ), .C(
        \Col_Fill[7][31] ), .D(\Col_Fill[7][30] ), .Q(n3030) );
  NOR40 U74228 ( .A(\Col_Fill[0][12] ), .B(\Col_Fill[0][11] ), .C(
        \Col_Fill[0][10] ), .D(\Col_Fill[0][0] ), .Q(n3076) );
  NOR40 U74229 ( .A(\Col_Fill[1][13] ), .B(\Col_Fill[1][12] ), .C(
        \Col_Fill[1][11] ), .D(\Col_Fill[1][10] ), .Q(n3087) );
  NOR40 U74230 ( .A(\Col_Fill[1][0] ), .B(\Col_Fill[0][9] ), .C(
        \Col_Fill[0][8] ), .D(\Col_Fill[0][7] ), .Q(n3086) );
  NOR40 U74231 ( .A(\Col_Fill[1][28] ), .B(\Col_Fill[1][27] ), .C(
        \Col_Fill[1][26] ), .D(\Col_Fill[1][25] ), .Q(n3091) );
  NOR40 U74232 ( .A(\Col_Fill[1][24] ), .B(\Col_Fill[1][23] ), .C(
        \Col_Fill[1][22] ), .D(\Col_Fill[1][21] ), .Q(n3090) );
  NOR40 U74233 ( .A(\Col_Fill[1][17] ), .B(\Col_Fill[1][16] ), .C(
        \Col_Fill[1][15] ), .D(\Col_Fill[1][14] ), .Q(n3088) );
  NOR40 U74234 ( .A(\Col_Fill[1][31] ), .B(\Col_Fill[1][30] ), .C(
        \Col_Fill[1][2] ), .D(\Col_Fill[1][29] ), .Q(n3092) );
  AOI311 U74235 ( .A(n65604), .B(n65577), .C(n65610), .D(n66580), .Q(N4434) );
  AOI311 U74236 ( .A(n65604), .B(N3200), .C(m[2]), .D(n66580), .Q(N4847) );
  BUF6 U74237 ( .A(n[5]), .Q(n65601) );
  OAI311 U74238 ( .A(n3476), .B(C4_OUT[1]), .C(C4_OUT[0]), .D(n3720), .Q(N2630) );
  NAND22 U74239 ( .A(start), .B(n3274), .Q(n3720) );
  NAND22 U74240 ( .A(n66685), .B(n66684), .Q(N3195) );
  AOI211 U74241 ( .A(n65604), .B(N3200), .C(n65610), .Q(n66685) );
  NOR21 U74242 ( .A(n1682), .B(C4_OUT[1]), .Q(n3655) );
  INV3 U74243 ( .A(N3200), .Q(n65584) );
  NOR21 U74244 ( .A(n1681), .B(C4_OUT[0]), .Q(n3676) );
  NOR21 U74245 ( .A(state[0]), .B(state[1]), .Q(n3274) );
  BUF2 U74246 ( .A(\OFill[23][0] ), .Q(n65651) );
  BUF2 U74247 ( .A(\OFill[21][0] ), .Q(n65649) );
  BUF2 U74248 ( .A(\OFill[7][0] ), .Q(n65667) );
  BUF2 U74249 ( .A(\OFill[5][0] ), .Q(n65665) );
  BUF2 U74250 ( .A(\OFill[55][0] ), .Q(n65619) );
  BUF2 U74251 ( .A(\OFill[53][0] ), .Q(n65617) );
  BUF2 U74252 ( .A(\OFill[39][0] ), .Q(n65635) );
  BUF2 U74253 ( .A(\OFill[37][0] ), .Q(n65633) );
  BUF2 U74254 ( .A(\GFill[23][0] ), .Q(n65715) );
  BUF2 U74255 ( .A(\GFill[21][0] ), .Q(n65713) );
  BUF2 U74256 ( .A(\GFill[7][0] ), .Q(n65731) );
  BUF2 U74257 ( .A(\GFill[5][0] ), .Q(n65729) );
  BUF2 U74258 ( .A(\GFill[55][0] ), .Q(n65683) );
  BUF2 U74259 ( .A(\GFill[53][0] ), .Q(n65681) );
  BUF2 U74260 ( .A(\GFill[39][0] ), .Q(n65699) );
  BUF2 U74261 ( .A(\GFill[37][0] ), .Q(n65697) );
  BUF2 U74262 ( .A(\OFill[19][0] ), .Q(n65647) );
  BUF2 U74263 ( .A(\OFill[17][0] ), .Q(n65645) );
  BUF2 U74264 ( .A(\OFill[31][0] ), .Q(n65659) );
  BUF2 U74265 ( .A(\OFill[29][0] ), .Q(n65657) );
  BUF2 U74266 ( .A(\OFill[27][0] ), .Q(n65655) );
  BUF2 U74267 ( .A(\OFill[25][0] ), .Q(n65653) );
  BUF2 U74268 ( .A(\OFill[3][0] ), .Q(n65663) );
  BUF2 U74269 ( .A(\OFill[1][0] ), .Q(n65661) );
  BUF2 U74270 ( .A(\OFill[15][0] ), .Q(n65675) );
  BUF2 U74271 ( .A(\OFill[13][0] ), .Q(n65673) );
  BUF2 U74272 ( .A(\OFill[11][0] ), .Q(n65671) );
  BUF2 U74273 ( .A(\OFill[9][0] ), .Q(n65669) );
  BUF2 U74274 ( .A(\OFill[51][0] ), .Q(n65615) );
  BUF2 U74275 ( .A(\OFill[49][0] ), .Q(n65613) );
  BUF2 U74276 ( .A(\OFill[63][0] ), .Q(n65627) );
  BUF2 U74277 ( .A(\OFill[61][0] ), .Q(n65625) );
  BUF2 U74278 ( .A(\OFill[59][0] ), .Q(n65623) );
  BUF2 U74279 ( .A(\OFill[57][0] ), .Q(n65621) );
  BUF2 U74280 ( .A(\OFill[35][0] ), .Q(n65631) );
  BUF2 U74281 ( .A(\OFill[33][0] ), .Q(n65629) );
  BUF2 U74282 ( .A(\OFill[47][0] ), .Q(n65643) );
  BUF2 U74283 ( .A(\OFill[45][0] ), .Q(n65641) );
  BUF2 U74284 ( .A(\OFill[43][0] ), .Q(n65639) );
  BUF2 U74285 ( .A(\OFill[41][0] ), .Q(n65637) );
  BUF2 U74286 ( .A(\GFill[19][0] ), .Q(n65711) );
  BUF2 U74287 ( .A(\GFill[17][0] ), .Q(n65709) );
  BUF2 U74288 ( .A(\GFill[31][0] ), .Q(n65723) );
  BUF2 U74289 ( .A(\GFill[29][0] ), .Q(n65721) );
  BUF2 U74290 ( .A(\GFill[27][0] ), .Q(n65719) );
  BUF2 U74291 ( .A(\GFill[25][0] ), .Q(n65717) );
  BUF2 U74292 ( .A(\GFill[3][0] ), .Q(n65727) );
  BUF2 U74293 ( .A(\GFill[1][0] ), .Q(n65725) );
  BUF2 U74294 ( .A(\GFill[15][0] ), .Q(n65739) );
  BUF2 U74295 ( .A(\GFill[13][0] ), .Q(n65737) );
  BUF2 U74296 ( .A(\GFill[11][0] ), .Q(n65735) );
  BUF2 U74297 ( .A(\GFill[9][0] ), .Q(n65733) );
  BUF2 U74298 ( .A(\GFill[51][0] ), .Q(n65679) );
  BUF2 U74299 ( .A(\GFill[49][0] ), .Q(n65677) );
  BUF2 U74300 ( .A(\GFill[63][0] ), .Q(n65691) );
  BUF2 U74301 ( .A(\GFill[61][0] ), .Q(n65689) );
  BUF2 U74302 ( .A(\GFill[59][0] ), .Q(n65687) );
  BUF2 U74303 ( .A(\GFill[57][0] ), .Q(n65685) );
  BUF2 U74304 ( .A(\GFill[35][0] ), .Q(n65695) );
  BUF2 U74305 ( .A(\GFill[33][0] ), .Q(n65693) );
  BUF2 U74306 ( .A(\GFill[47][0] ), .Q(n65707) );
  BUF2 U74307 ( .A(\GFill[45][0] ), .Q(n65705) );
  BUF2 U74308 ( .A(\GFill[43][0] ), .Q(n65703) );
  BUF2 U74309 ( .A(\GFill[41][0] ), .Q(n65701) );
  NOR21 U74310 ( .A(n3079), .B(n3080), .Q(n3078) );
  NAND41 U74311 ( .A(\Col_Fill[7][3] ), .B(\Col_Fill[6][3] ), .C(
        \Col_Fill[5][3] ), .D(\Col_Fill[4][3] ), .Q(n3080) );
  NAND41 U74312 ( .A(\Col_Fill[3][3] ), .B(\Col_Fill[2][3] ), .C(
        \Col_Fill[1][3] ), .D(\Col_Fill[0][3] ), .Q(n3079) );
  INV3 U74313 ( .A(N3200), .Q(n65585) );
  BUF2 U74314 ( .A(\OFill[20][0] ), .Q(n65648) );
  BUF2 U74315 ( .A(\OFill[16][0] ), .Q(n65644) );
  BUF2 U74316 ( .A(\OFill[28][0] ), .Q(n65656) );
  BUF2 U74317 ( .A(\OFill[24][0] ), .Q(n65652) );
  BUF2 U74318 ( .A(\OFill[4][0] ), .Q(n65664) );
  BUF2 U74319 ( .A(\OFill[0][0] ), .Q(n65660) );
  BUF2 U74320 ( .A(\OFill[12][0] ), .Q(n65672) );
  BUF2 U74321 ( .A(\OFill[8][0] ), .Q(n65668) );
  BUF2 U74322 ( .A(\OFill[52][0] ), .Q(n65616) );
  BUF2 U74323 ( .A(\OFill[48][0] ), .Q(n65612) );
  BUF2 U74324 ( .A(\OFill[60][0] ), .Q(n65624) );
  BUF2 U74325 ( .A(\OFill[56][0] ), .Q(n65620) );
  BUF2 U74326 ( .A(\OFill[36][0] ), .Q(n65632) );
  BUF2 U74327 ( .A(\OFill[32][0] ), .Q(n65628) );
  BUF2 U74328 ( .A(\OFill[44][0] ), .Q(n65640) );
  BUF2 U74329 ( .A(\OFill[40][0] ), .Q(n65636) );
  BUF2 U74330 ( .A(\GFill[20][0] ), .Q(n65712) );
  BUF2 U74331 ( .A(\GFill[16][0] ), .Q(n65708) );
  BUF2 U74332 ( .A(\GFill[28][0] ), .Q(n65720) );
  BUF2 U74333 ( .A(\GFill[24][0] ), .Q(n65716) );
  BUF2 U74334 ( .A(\GFill[4][0] ), .Q(n65728) );
  BUF2 U74335 ( .A(\GFill[0][0] ), .Q(n65724) );
  BUF2 U74336 ( .A(\GFill[12][0] ), .Q(n65736) );
  BUF2 U74337 ( .A(\GFill[8][0] ), .Q(n65732) );
  BUF2 U74338 ( .A(\GFill[52][0] ), .Q(n65680) );
  BUF2 U74339 ( .A(\GFill[48][0] ), .Q(n65676) );
  BUF2 U74340 ( .A(\GFill[60][0] ), .Q(n65688) );
  BUF2 U74341 ( .A(\GFill[56][0] ), .Q(n65684) );
  BUF2 U74342 ( .A(\GFill[36][0] ), .Q(n65696) );
  BUF2 U74343 ( .A(\GFill[32][0] ), .Q(n65692) );
  BUF2 U74344 ( .A(\GFill[44][0] ), .Q(n65704) );
  BUF2 U74345 ( .A(\GFill[40][0] ), .Q(n65700) );
  INV3 U74346 ( .A(N1208), .Q(n65781) );
  INV3 U74347 ( .A(N1167), .Q(n65920) );
  INV3 U74348 ( .A(m[1]), .Q(n65608) );
  INV3 U74349 ( .A(n[3]), .Q(n65596) );
  INV3 U74350 ( .A(m[2]), .Q(n65611) );
  LOGIC0 U74351 ( .Q(n65544) );
  LOGIC1 U74352 ( .Q(n807) );
  OAI212 U74353 ( .A(n65829), .B(n65770), .C(n66097), .Q(N740) );
  OAI212 U74354 ( .A(n65818), .B(n65774), .C(n66097), .Q(N1010) );
  OAI212 U74355 ( .A(n65789), .B(n65780), .C(n66114), .Q(N1004) );
  OAI212 U74356 ( .A(n65831), .B(n65759), .C(n66103), .Q(N722) );
  OAI212 U74357 ( .A(n65784), .B(n65771), .C(n66097), .Q(N716) );
  OAI212 U74358 ( .A(n65782), .B(n65774), .C(n66114), .Q(N980) );
  OAI212 U74359 ( .A(n65807), .B(n65777), .C(n66114), .Q(N704) );
  CLKIN3 U74360 ( .A(n65885), .Q(n65782) );
  CLKIN3 U74361 ( .A(n65910), .Q(n65783) );
  CLKIN3 U74362 ( .A(n65855), .Q(n65784) );
  CLKIN3 U74363 ( .A(n65869), .Q(n65785) );
  CLKIN3 U74364 ( .A(n65840), .Q(n65786) );
  CLKIN3 U74365 ( .A(n65839), .Q(n65787) );
  CLKIN3 U74366 ( .A(n65901), .Q(n65788) );
  CLKIN3 U74367 ( .A(n65843), .Q(n65789) );
  CLKIN3 U74368 ( .A(n65903), .Q(n65790) );
  CLKIN3 U74369 ( .A(n65899), .Q(n65791) );
  CLKIN3 U74370 ( .A(n65874), .Q(n65792) );
  CLKIN3 U74371 ( .A(n65873), .Q(n65793) );
  CLKIN3 U74372 ( .A(n65862), .Q(n65794) );
  CLKIN3 U74373 ( .A(n65852), .Q(n65795) );
  CLKIN3 U74374 ( .A(n65872), .Q(n65796) );
  CLKIN3 U74375 ( .A(n65846), .Q(n65797) );
  CLKIN3 U74376 ( .A(n65844), .Q(n65798) );
  CLKIN3 U74377 ( .A(n65846), .Q(n65799) );
  CLKIN3 U74378 ( .A(n65851), .Q(n65800) );
  CLKIN3 U74379 ( .A(n65848), .Q(n65801) );
  CLKIN3 U74380 ( .A(n65845), .Q(n65802) );
  CLKIN3 U74381 ( .A(n65850), .Q(n65803) );
  CLKIN3 U74382 ( .A(n65847), .Q(n65804) );
  CLKIN3 U74383 ( .A(n65852), .Q(n65805) );
  CLKIN3 U74384 ( .A(n65849), .Q(n65806) );
  CLKIN3 U74385 ( .A(n65856), .Q(n65807) );
  CLKIN3 U74386 ( .A(n65906), .Q(n65808) );
  CLKIN3 U74387 ( .A(n65865), .Q(n65809) );
  CLKIN3 U74388 ( .A(n65857), .Q(n65810) );
  CLKIN3 U74389 ( .A(n65858), .Q(n65811) );
  CLKIN3 U74390 ( .A(n65860), .Q(n65812) );
  CLKIN3 U74391 ( .A(n65861), .Q(n65813) );
  CLKIN3 U74392 ( .A(n65862), .Q(n65814) );
  CLKIN3 U74393 ( .A(n65863), .Q(n65815) );
  CLKIN3 U74394 ( .A(n65864), .Q(n65816) );
  CLKIN3 U74395 ( .A(n65865), .Q(n65817) );
  CLKIN3 U74396 ( .A(n65866), .Q(n65818) );
  CLKIN3 U74397 ( .A(n65867), .Q(n65819) );
  CLKIN3 U74398 ( .A(n65868), .Q(n65820) );
  CLKIN3 U74399 ( .A(n65843), .Q(n65821) );
  CLKIN3 U74400 ( .A(n65902), .Q(n65822) );
  CLKIN3 U74401 ( .A(n65855), .Q(n65823) );
  CLKIN3 U74402 ( .A(n65862), .Q(n65824) );
  CLKIN3 U74403 ( .A(n65854), .Q(n65825) );
  CLKIN3 U74404 ( .A(n65871), .Q(n65826) );
  CLKIN3 U74405 ( .A(n65908), .Q(n65827) );
  CLKIN3 U74406 ( .A(n65871), .Q(n65828) );
  CLKIN3 U74407 ( .A(n65870), .Q(n65829) );
  CLKIN3 U74408 ( .A(n65897), .Q(n65830) );
  CLKIN3 U74409 ( .A(n65869), .Q(n65831) );
  XOR20 U74410 ( .A(n65963), .B(\sub_140_2_cf/carry [10]), .Q(N1524) );
  NAND20 U74411 ( .A(n65963), .B(\sub_140_2_cf/carry [9]), .Q(n65956) );
  XOR20 U74412 ( .A(n65963), .B(\sub_140_2_cf/carry [9]), .Q(N1523) );
  CLKIN0 U74413 ( .A(n65956), .Q(\sub_140_2_cf/carry [10]) );
  NAND20 U74414 ( .A(n65963), .B(\sub_140_2_cf/carry [8]), .Q(n65957) );
  XOR20 U74415 ( .A(n65963), .B(\sub_140_2_cf/carry [8]), .Q(N1522) );
  CLKIN0 U74416 ( .A(n65957), .Q(\sub_140_2_cf/carry [9]) );
  NAND20 U74417 ( .A(n65963), .B(\sub_140_2_cf/carry [7]), .Q(n65958) );
  XOR20 U74418 ( .A(n65963), .B(\sub_140_2_cf/carry [7]), .Q(N1521) );
  CLKIN0 U74419 ( .A(n65958), .Q(\sub_140_2_cf/carry [8]) );
  NAND20 U74420 ( .A(n65963), .B(\sub_140_2_cf/carry [6]), .Q(n65959) );
  XOR20 U74421 ( .A(n65963), .B(\sub_140_2_cf/carry [6]), .Q(N1520) );
  CLKIN0 U74422 ( .A(n65959), .Q(\sub_140_2_cf/carry [7]) );
  NAND20 U74423 ( .A(N11202), .B(\sub_140_2_cf/carry [5]), .Q(n65960) );
  XOR20 U74424 ( .A(N11202), .B(\sub_140_2_cf/carry [5]), .Q(N1519) );
  CLKIN0 U74425 ( .A(n65960), .Q(\sub_140_2_cf/carry [6]) );
  NOR20 U74426 ( .A(\sub_140_2_cf/carry [4]), .B(N11203), .Q(n65961) );
  XNR20 U74427 ( .A(\sub_140_2_cf/carry [4]), .B(N11203), .Q(N1518) );
  CLKIN0 U74428 ( .A(n65961), .Q(\sub_140_2_cf/carry [5]) );
  NOR20 U74429 ( .A(\sub_140_2_cf/carry [3]), .B(N11204), .Q(n65962) );
  XNR20 U74430 ( .A(\sub_140_2_cf/carry [3]), .B(N11204), .Q(N1517) );
  CLKIN0 U74431 ( .A(n65962), .Q(\sub_140_2_cf/carry [4]) );
  XOR20 U74432 ( .A(n66108), .B(\sub_140_b0/carry [5]), .Q(N11202) );
  NAND20 U74433 ( .A(n66107), .B(\sub_140_b0/carry [4]), .Q(n65964) );
  XOR20 U74434 ( .A(n66107), .B(\sub_140_b0/carry [4]), .Q(N11203) );
  CLKIN0 U74435 ( .A(n65964), .Q(\sub_140_b0/carry [5]) );
  NAND20 U74436 ( .A(n66106), .B(\sub_140_b0/carry [3]), .Q(n65965) );
  XOR20 U74437 ( .A(n66106), .B(\sub_140_b0/carry [3]), .Q(N11204) );
  CLKIN0 U74438 ( .A(n65965), .Q(\sub_140_b0/carry [4]) );
  NAND20 U74439 ( .A(N11205), .B(N11206), .Q(n65966) );
  XOR20 U74440 ( .A(N11205), .B(N11206), .Q(N1516) );
  CLKIN0 U74441 ( .A(n65966), .Q(\sub_140_2_cf/carry [3]) );
  NAND20 U74442 ( .A(n66105), .B(\sub_140_b0/carry [2]), .Q(n65967) );
  XOR20 U74443 ( .A(n66105), .B(\sub_140_b0/carry [2]), .Q(N11205) );
  CLKIN0 U74444 ( .A(n65967), .Q(\sub_140_b0/carry [3]) );
  NAND20 U74445 ( .A(n66104), .B(n65420), .Q(n65968) );
  CLKIN0 U74446 ( .A(n65968), .Q(\sub_140_b0/carry [2]) );
  XOR20 U74447 ( .A(n65976), .B(\sub_171_2_cf/carry[10] ), .Q(N2067) );
  NAND20 U74448 ( .A(n65976), .B(\sub_171_2_cf/carry[9] ), .Q(n65969) );
  XOR20 U74449 ( .A(n65976), .B(\sub_171_2_cf/carry[9] ), .Q(N2066) );
  CLKIN0 U74450 ( .A(n65969), .Q(\sub_171_2_cf/carry[10] ) );
  NAND20 U74451 ( .A(n65976), .B(\sub_171_2_cf/carry[8] ), .Q(n65970) );
  XOR20 U74452 ( .A(n65976), .B(\sub_171_2_cf/carry[8] ), .Q(N2065) );
  CLKIN0 U74453 ( .A(n65970), .Q(\sub_171_2_cf/carry[9] ) );
  NAND20 U74454 ( .A(n65976), .B(\sub_171_2_cf/carry[7] ), .Q(n65971) );
  XOR20 U74455 ( .A(n65976), .B(\sub_171_2_cf/carry[7] ), .Q(N2064) );
  CLKIN0 U74456 ( .A(n65971), .Q(\sub_171_2_cf/carry[8] ) );
  NAND20 U74457 ( .A(n65976), .B(\sub_171_2_cf/carry[6] ), .Q(n65972) );
  XOR20 U74458 ( .A(n65976), .B(\sub_171_2_cf/carry[6] ), .Q(N2063) );
  CLKIN0 U74459 ( .A(n65972), .Q(\sub_171_2_cf/carry[7] ) );
  NAND20 U74460 ( .A(N11212), .B(\sub_171_2_cf/carry[5] ), .Q(n65973) );
  XOR20 U74461 ( .A(N11212), .B(\sub_171_2_cf/carry[5] ), .Q(N2062) );
  CLKIN0 U74462 ( .A(n65973), .Q(\sub_171_2_cf/carry[6] ) );
  NOR20 U74463 ( .A(\sub_171_2_cf/carry[4] ), .B(N11213), .Q(n65974) );
  XNR20 U74464 ( .A(\sub_171_2_cf/carry[4] ), .B(N11213), .Q(N2061) );
  CLKIN0 U74465 ( .A(n65974), .Q(\sub_171_2_cf/carry[5] ) );
  NOR20 U74466 ( .A(\sub_171_2_cf/carry[3] ), .B(N11214), .Q(n65975) );
  XNR20 U74467 ( .A(\sub_171_2_cf/carry[3] ), .B(N11214), .Q(N2060) );
  CLKIN0 U74468 ( .A(n65975), .Q(\sub_171_2_cf/carry[4] ) );
  XOR20 U74469 ( .A(n66122), .B(\sub_171_b0/carry [5]), .Q(N11212) );
  NAND20 U74470 ( .A(n66121), .B(\sub_171_b0/carry [4]), .Q(n65977) );
  XOR20 U74471 ( .A(n66121), .B(\sub_171_b0/carry [4]), .Q(N11213) );
  CLKIN0 U74472 ( .A(n65977), .Q(\sub_171_b0/carry [5]) );
  NAND20 U74473 ( .A(n66120), .B(\sub_171_b0/carry [3]), .Q(n65978) );
  XOR20 U74474 ( .A(n66120), .B(\sub_171_b0/carry [3]), .Q(N11214) );
  CLKIN0 U74475 ( .A(n65978), .Q(\sub_171_b0/carry [4]) );
  NAND20 U74476 ( .A(N11215), .B(\sub_171_2_cf/carry[2] ), .Q(n65979) );
  XOR20 U74477 ( .A(N11215), .B(\sub_171_2_cf/carry[2] ), .Q(N2059) );
  CLKIN0 U74478 ( .A(n65979), .Q(\sub_171_2_cf/carry[3] ) );
  NAND20 U74479 ( .A(N11216), .B(n65740), .Q(n65980) );
  XOR20 U74480 ( .A(N11216), .B(n65740), .Q(N2058) );
  CLKIN0 U74481 ( .A(n65980), .Q(\sub_171_2_cf/carry[2] ) );
  NAND20 U74482 ( .A(n66119), .B(\sub_171_b0/carry [2]), .Q(n65981) );
  XOR20 U74483 ( .A(n66119), .B(\sub_171_b0/carry [2]), .Q(N11215) );
  CLKIN0 U74484 ( .A(n65981), .Q(\sub_171_b0/carry [3]) );
  NAND20 U74485 ( .A(n65451), .B(n65515), .Q(n65982) );
  XOR20 U74486 ( .A(n65451), .B(n65419), .Q(N11216) );
  CLKIN0 U74487 ( .A(n65982), .Q(\sub_171_b0/carry [2]) );
  XOR20 U74488 ( .A(n[3]), .B(n65580), .Q(N11520) );
  XOR20 U74489 ( .A(n[3]), .B(n65585), .Q(N11538) );
  XOR20 U74490 ( .A(n65601), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [5]), 
        .Q(N11542) );
  NAND20 U74491 ( .A(n[4]), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [4]), 
        .Q(n65983) );
  XOR20 U74492 ( .A(n65599), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [4]), 
        .Q(N11543) );
  CLKIN0 U74493 ( .A(n65983), .Q(\add_1_root_add_0_root_sub_348_9_cf/carry [5]) );
  NAND20 U74494 ( .A(N11544), .B(n65579), .Q(n65984) );
  CLKIN0 U74495 ( .A(n65984), .Q(\add_0_root_add_0_root_sub_348_9_cf/carry [4]) );
  NAND20 U74496 ( .A(n[3]), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [3]), 
        .Q(n65985) );
  XOR20 U74497 ( .A(n[3]), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [3]), 
        .Q(N11544) );
  NAND20 U74498 ( .A(n65916), .B(n65746), .Q(n65986) );
  XNR20 U74499 ( .A(n65601), .B(\r11553/carry[5] ), .Q(N11404) );
  XNR20 U74500 ( .A(\add_1_root_add_0_root_sub_331_4_cf/carry[4] ), .B(n65599), 
        .Q(N11405) );
  NAND20 U74501 ( .A(N11406), .B(n65579), .Q(n65987) );
  CLKIN0 U74502 ( .A(n65987), .Q(\add_0_root_add_0_root_sub_331_4_cf/carry [4]) );
  NOR20 U74503 ( .A(\r34786/carry [3]), .B(n65594), .Q(n65988) );
  XNR20 U74504 ( .A(\r34786/carry [3]), .B(n[3]), .Q(N11406) );
  XNR20 U74505 ( .A(n65601), .B(\r34786/carry [5]), .Q(N11380) );
  XNR20 U74506 ( .A(\add_1_root_add_0_root_sub_328_4_cf/carry[4] ), .B(n65599), 
        .Q(N11381) );
  NAND20 U74507 ( .A(N11382), .B(n65579), .Q(n65989) );
  CLKIN0 U74508 ( .A(n65989), .Q(\add_0_root_add_0_root_sub_328_4_cf/carry [4]) );
  NOR20 U74509 ( .A(\r34786/carry [3]), .B(n65594), .Q(n65990) );
  XNR20 U74510 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11382) );
  XNR20 U74511 ( .A(n65601), .B(\add_1_root_add_0_root_sub_328_8_cf/carry[5] ), 
        .Q(N11386) );
  NOR20 U74512 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[4] ), .B(n[4]), 
        .Q(n65991) );
  XNR20 U74513 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[4] ), .B(n65598), 
        .Q(N11387) );
  CLKIN0 U74514 ( .A(n65991), .Q(\add_1_root_add_0_root_sub_328_8_cf/carry[5] ) );
  NAND20 U74515 ( .A(N11388), .B(n65583), .Q(n65992) );
  CLKIN0 U74516 ( .A(n65992), .Q(\add_0_root_add_0_root_sub_328_8_cf/carry [4]) );
  XNR20 U74517 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[3] ), .B(n65593), 
        .Q(N11388) );
  NAND20 U74518 ( .A(n65744), .B(n65875), .Q(n65993) );
  XNR20 U74519 ( .A(N4042), .B(\add_1_root_add_0_root_sub_325_8_cf/carry[5] ), 
        .Q(N11356) );
  NOR20 U74520 ( .A(n65583), .B(N4041), .Q(n65994) );
  XNR20 U74521 ( .A(n65580), .B(N4041), .Q(N11357) );
  CLKIN0 U74522 ( .A(n65994), .Q(\add_1_root_add_0_root_sub_325_8_cf/carry[5] ) );
  NOR20 U74523 ( .A(N1167), .B(\add_0_root_add_0_root_sub_325_8_cf/carry [2]), 
        .Q(n65995) );
  CLKIN0 U74524 ( .A(n65995), .Q(\add_0_root_add_0_root_sub_325_8_cf/carry [3]) );
  NAND20 U74525 ( .A(n65906), .B(n65745), .Q(n65996) );
  CLKIN0 U74526 ( .A(n65996), .Q(\add_0_root_add_0_root_sub_325_8_cf/carry [2]) );
  XNR20 U74527 ( .A(n65611), .B(\add_1_root_add_0_root_sub_325_12_cf/carry[5] ), .Q(N11362) );
  NOR20 U74528 ( .A(n65578), .B(n65604), .Q(n65997) );
  XNR20 U74529 ( .A(n65578), .B(n65604), .Q(N11363) );
  CLKIN0 U74530 ( .A(n65997), .Q(
        \add_1_root_add_0_root_sub_325_12_cf/carry[5] ) );
  XNR20 U74531 ( .A(N4030), .B(\add_1_root_add_0_root_sub_325_4_cf/carry[5] ), 
        .Q(N11350) );
  NOR20 U74532 ( .A(n65578), .B(n65607), .Q(n65998) );
  XNR20 U74533 ( .A(n65578), .B(n65606), .Q(N11351) );
  CLKIN0 U74534 ( .A(n65998), .Q(\add_1_root_add_0_root_sub_325_4_cf/carry[5] ) );
  NOR20 U74535 ( .A(N1167), .B(N1208), .Q(n65999) );
  CLKIN0 U74536 ( .A(n65999), .Q(\add_0_root_add_0_root_sub_325_4_cf/carry [3]) );
  NOR20 U74537 ( .A(N1167), .B(n66114), .Q(n66000) );
  CLKIN0 U74538 ( .A(n66000), .Q(\add_0_root_sub_0_root_sub_297_3/carry [3])
         );
  NOR20 U74539 ( .A(N1167), .B(n66097), .Q(n66001) );
  CLKIN0 U74540 ( .A(n66001), .Q(\add_0_root_sub_0_root_sub_297_6/carry [3])
         );
  NAND20 U74541 ( .A(N2936), .B(n65579), .Q(n66002) );
  CLKIN0 U74542 ( .A(n66002), .Q(\add_0_root_sub_0_root_sub_297_9/carry [4])
         );
  NAND20 U74543 ( .A(N3072), .B(n65579), .Q(n66003) );
  CLKIN0 U74544 ( .A(n66003), .Q(\add_0_root_sub_0_root_sub_300_5/carry [4])
         );
  NAND20 U74545 ( .A(N3090), .B(n65581), .Q(n66004) );
  CLKIN0 U74546 ( .A(n66004), .Q(\add_0_root_sub_0_root_sub_300_8/carry [4])
         );
  NAND20 U74547 ( .A(N3245), .B(n65579), .Q(n66005) );
  CLKIN0 U74548 ( .A(n66005), .Q(\add_0_root_sub_0_root_sub_303_7/carry [4])
         );
  XOR20 U74549 ( .A(n65601), .B(\r40165/carry[5] ), .Q(N11434) );
  NAND20 U74550 ( .A(n[4]), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [4]), 
        .Q(n66006) );
  XOR20 U74551 ( .A(n65599), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [4]), 
        .Q(N11435) );
  CLKIN0 U74552 ( .A(n66006), .Q(\r40165/carry[5] ) );
  NAND20 U74553 ( .A(N11436), .B(n65579), .Q(n66007) );
  CLKIN0 U74554 ( .A(n66007), .Q(\r40166/carry [4]) );
  XOR20 U74555 ( .A(n[3]), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [3]), 
        .Q(N11436) );
  NAND20 U74556 ( .A(n[3]), .B(n65585), .Q(n66008) );
  XOR20 U74557 ( .A(n65594), .B(n65584), .Q(N11430) );
  XNR20 U74558 ( .A(n65601), .B(\r11555/carry[5] ), .Q(N11470) );
  XNR20 U74559 ( .A(\r41369/carry[4] ), .B(n65599), .Q(N11471) );
  NAND20 U74560 ( .A(N11472), .B(n65579), .Q(n66009) );
  CLKIN0 U74561 ( .A(n66009), .Q(\r41370/carry [4]) );
  NOR20 U74562 ( .A(N1167), .B(n65594), .Q(n66010) );
  XNR20 U74563 ( .A(n65915), .B(n65593), .Q(N11472) );
  XNR20 U74564 ( .A(n65601), .B(\add_1_root_add_0_root_sub_403_4_cf/carry[5] ), 
        .Q(N11458) );
  XNR20 U74565 ( .A(\add_1_root_add_0_root_sub_331_4_cf/carry[4] ), .B(n65599), 
        .Q(N11459) );
  NAND20 U74566 ( .A(N11460), .B(n65579), .Q(n66011) );
  CLKIN0 U74567 ( .A(n66011), .Q(\r38962/carry [4]) );
  XNR20 U74568 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11460) );
  XNR20 U74569 ( .A(n65601), .B(\r30598/carry[5] ), .Q(N11464) );
  NOR20 U74570 ( .A(\r30598/carry[4] ), .B(n[4]), .Q(n66012) );
  XNR20 U74571 ( .A(\r30598/carry[4] ), .B(n65598), .Q(N11465) );
  CLKIN0 U74572 ( .A(n66012), .Q(\r30598/carry[5] ) );
  NAND20 U74573 ( .A(N11466), .B(n65580), .Q(n66013) );
  CLKIN0 U74574 ( .A(n66013), .Q(\r30599/carry [4]) );
  NOR20 U74575 ( .A(\r30598/carry[3] ), .B(n65594), .Q(n66014) );
  XNR20 U74576 ( .A(\r30598/carry[3] ), .B(n65594), .Q(N11466) );
  CLKIN0 U74577 ( .A(n66014), .Q(\r30598/carry[4] ) );
  NOR20 U74578 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65915), 
        .Q(n66015) );
  CLKIN0 U74579 ( .A(n66015), .Q(\r30598/carry[3] ) );
  XNR20 U74580 ( .A(n65601), .B(\r34786/carry [5]), .Q(N11488) );
  NOR20 U74581 ( .A(\add_1_root_add_0_root_sub_328_4_cf/carry[4] ), .B(n[4]), 
        .Q(n66016) );
  XNR20 U74582 ( .A(\add_1_root_add_0_root_sub_328_4_cf/carry[4] ), .B(n65599), 
        .Q(N11489) );
  CLKIN0 U74583 ( .A(n66016), .Q(\r34786/carry [5]) );
  NAND20 U74584 ( .A(N11490), .B(n65578), .Q(n66017) );
  CLKIN0 U74585 ( .A(n66017), .Q(\r34787/carry [4]) );
  XNR20 U74586 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11490) );
  NOR20 U74587 ( .A(n65757), .B(n65915), .Q(n66018) );
  XNR20 U74588 ( .A(n65601), .B(\r33598/carry[5] ), .Q(N11494) );
  NOR20 U74589 ( .A(\r33598/carry[4] ), .B(n65599), .Q(n66019) );
  XNR20 U74590 ( .A(\r33598/carry[4] ), .B(n65598), .Q(N11495) );
  CLKIN0 U74591 ( .A(n66019), .Q(\r33598/carry[5] ) );
  NAND20 U74592 ( .A(N11496), .B(n65584), .Q(n66020) );
  CLKIN0 U74593 ( .A(n66020), .Q(\r33599/carry [4]) );
  NOR20 U74594 ( .A(\r30598/carry[3] ), .B(n65594), .Q(n66021) );
  XNR20 U74595 ( .A(\r12189/carry[3] ), .B(n65594), .Q(N11496) );
  CLKIN0 U74596 ( .A(n66021), .Q(\r33598/carry[4] ) );
  XOR20 U74597 ( .A(n65758), .B(n65844), .Q(N1220) );
  XOR20 U74598 ( .A(n65601), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [5]), 
        .Q(N11530) );
  XOR20 U74599 ( .A(n65599), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [4]), 
        .Q(N11531) );
  NAND20 U74600 ( .A(N11532), .B(n65578), .Q(n66022) );
  CLKIN0 U74601 ( .A(n66022), .Q(\add_0_root_add_0_root_sub_420_9_cf/carry [4]) );
  XOR20 U74602 ( .A(n65594), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [3]), 
        .Q(N11532) );
  XOR20 U74603 ( .A(n65916), .B(n65758), .Q(N1263) );
  XOR20 U74604 ( .A(n65594), .B(n65582), .Q(N11526) );
  XOR20 U74605 ( .A(n65594), .B(n65580), .Q(N11508) );
  XNR20 U74606 ( .A(n65601), .B(\r39563/carry[5] ), .Q(N11512) );
  NOR20 U74607 ( .A(\add_1_root_add_0_root_sub_328_4_cf/carry[4] ), .B(n[4]), 
        .Q(n66023) );
  XNR20 U74608 ( .A(\add_1_root_add_0_root_sub_331_4_cf/carry[4] ), .B(n65599), 
        .Q(N11513) );
  CLKIN0 U74609 ( .A(n66023), .Q(\r39563/carry[5] ) );
  NAND20 U74610 ( .A(N11514), .B(n65578), .Q(n66024) );
  CLKIN0 U74611 ( .A(n66024), .Q(\r39564/carry [4]) );
  XNR20 U74612 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11514) );
  XNR20 U74613 ( .A(n65601), .B(\add_1_root_add_0_root_sub_403_4_cf/carry[5] ), 
        .Q(N11392) );
  NOR20 U74614 ( .A(\add_1_root_add_0_root_sub_331_4_cf/carry[4] ), .B(n65599), 
        .Q(n66025) );
  XNR20 U74615 ( .A(\r12188/carry [4]), .B(n65598), .Q(N11393) );
  CLKIN0 U74616 ( .A(n66025), .Q(\add_1_root_add_0_root_sub_403_4_cf/carry[5] ) );
  NAND20 U74617 ( .A(N11394), .B(n65578), .Q(n66026) );
  CLKIN0 U74618 ( .A(n66026), .Q(\add_0_root_add_0_root_sub_403_4_cf/carry [4]) );
  XNR20 U74619 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11394) );
  NAND20 U74620 ( .A(n[3]), .B(n65578), .Q(n66027) );
  XNR20 U74621 ( .A(n65601), .B(\add_1_root_add_0_root_sub_400_4_cf/carry[5] ), 
        .Q(N11368) );
  NOR20 U74622 ( .A(\add_1_root_add_0_root_sub_331_4_cf/carry[4] ), .B(n65599), 
        .Q(n66028) );
  XNR20 U74623 ( .A(\add_1_root_add_0_root_sub_328_4_cf/carry[4] ), .B(n65599), 
        .Q(N11369) );
  CLKIN0 U74624 ( .A(n66028), .Q(\add_1_root_add_0_root_sub_400_4_cf/carry[5] ) );
  NAND20 U74625 ( .A(N11370), .B(n65578), .Q(n66029) );
  CLKIN0 U74626 ( .A(n66029), .Q(\add_0_root_add_0_root_sub_400_4_cf/carry [4]) );
  XNR20 U74627 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11370) );
  XNR20 U74628 ( .A(n65601), .B(\add_1_root_add_0_root_sub_400_8_cf/carry[5] ), 
        .Q(N11374) );
  NOR20 U74629 ( .A(\r12189/carry[4] ), .B(n[4]), .Q(n66030) );
  XNR20 U74630 ( .A(\r12189/carry[4] ), .B(n65598), .Q(N11375) );
  CLKIN0 U74631 ( .A(n66030), .Q(\add_1_root_add_0_root_sub_400_8_cf/carry[5] ) );
  NAND20 U74632 ( .A(N11376), .B(n65581), .Q(n66031) );
  CLKIN0 U74633 ( .A(n66031), .Q(\add_0_root_add_0_root_sub_400_8_cf/carry [4]) );
  XNR20 U74634 ( .A(\r30598/carry[3] ), .B(n65594), .Q(N11376) );
  XNR20 U74635 ( .A(n65601), .B(\r11555/carry[5] ), .Q(N11344) );
  XNR20 U74636 ( .A(\r41369/carry[4] ), .B(n65598), .Q(N11345) );
  NAND20 U74637 ( .A(N11346), .B(n65578), .Q(n66032) );
  CLKIN0 U74638 ( .A(n66032), .Q(
        \add_0_root_add_0_root_sub_397_12_cf/carry [4]) );
  XNR20 U74639 ( .A(N1167), .B(n65594), .Q(N11346) );
  XNR20 U74640 ( .A(n65601), .B(\add_1_root_add_0_root_sub_403_4_cf/carry[5] ), 
        .Q(N11332) );
  XNR20 U74641 ( .A(\r12188/carry [4]), .B(n65599), .Q(N11333) );
  NAND20 U74642 ( .A(N11334), .B(n65578), .Q(n66033) );
  CLKIN0 U74643 ( .A(n66033), .Q(\add_0_root_add_0_root_sub_397_4_cf/carry [4]) );
  XNR20 U74644 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11334) );
  XNR20 U74645 ( .A(n65601), .B(\add_1_root_add_0_root_sub_328_8_cf/carry[5] ), 
        .Q(N11338) );
  XNR20 U74646 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[4] ), .B(n65598), 
        .Q(N11339) );
  NAND20 U74647 ( .A(N11340), .B(n65582), .Q(n66034) );
  CLKIN0 U74648 ( .A(n66034), .Q(\add_0_root_add_0_root_sub_397_8_cf/carry [4]) );
  NOR20 U74649 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[3] ), .B(n65594), 
        .Q(n66035) );
  XNR20 U74650 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[3] ), .B(n65594), 
        .Q(N11340) );
  NOR20 U74651 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(n65918), 
        .Q(n66036) );
  CLKIN0 U74652 ( .A(n66036), .Q(\add_1_root_add_0_root_sub_397_8_cf/carry[3] ) );
  XOR20 U74653 ( .A(n65601), .B(\r13448/carry[5] ), .Q(N11320) );
  NAND20 U74654 ( .A(n[4]), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [4]), 
        .Q(n66037) );
  XOR20 U74655 ( .A(n65598), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [4]), 
        .Q(N11321) );
  CLKIN0 U74656 ( .A(n66037), .Q(\r13448/carry[5] ) );
  NAND20 U74657 ( .A(N11322), .B(n65580), .Q(n66038) );
  CLKIN0 U74658 ( .A(n66038), .Q(\r13450/carry [4]) );
  XOR20 U74659 ( .A(n65594), .B(\add_1_root_add_0_root_sub_348_9_cf/carry [3]), 
        .Q(N11322) );
  XNR20 U74660 ( .A(n65601), .B(\r11555/carry[5] ), .Q(N11266) );
  NOR20 U74661 ( .A(\r41369/carry[4] ), .B(n65599), .Q(n66039) );
  XNR20 U74662 ( .A(\r41369/carry[4] ), .B(n65598), .Q(N11267) );
  CLKIN0 U74663 ( .A(n66039), .Q(\r11555/carry[5] ) );
  NAND20 U74664 ( .A(N11268), .B(n65580), .Q(n66040) );
  CLKIN0 U74665 ( .A(n66040), .Q(\r11558/carry [4]) );
  XNR20 U74666 ( .A(n65917), .B(n65594), .Q(N11268) );
  XNR20 U74667 ( .A(n65601), .B(\r11553/carry[5] ), .Q(N11254) );
  NOR20 U74668 ( .A(\add_1_root_add_0_root_sub_331_4_cf/carry[4] ), .B(n[4]), 
        .Q(n66041) );
  XNR20 U74669 ( .A(\r12188/carry [4]), .B(n65598), .Q(N11255) );
  CLKIN0 U74670 ( .A(n66041), .Q(\r11553/carry[5] ) );
  NAND20 U74671 ( .A(N11256), .B(n65584), .Q(n66042) );
  CLKIN0 U74672 ( .A(n66042), .Q(\r11556/carry [4]) );
  XNR20 U74673 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11256) );
  XNR20 U74674 ( .A(n65601), .B(\r11554/carry[5] ), .Q(N11260) );
  NOR20 U74675 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[4] ), .B(n[4]), 
        .Q(n66043) );
  XNR20 U74676 ( .A(\add_1_root_add_0_root_sub_397_8_cf/carry[4] ), .B(n65598), 
        .Q(N11261) );
  CLKIN0 U74677 ( .A(n66043), .Q(\r11554/carry[5] ) );
  NAND20 U74678 ( .A(N11262), .B(n65585), .Q(n66044) );
  CLKIN0 U74679 ( .A(n66044), .Q(\r11557/carry [4]) );
  XNR20 U74680 ( .A(\r12189/carry[3] ), .B(n65594), .Q(N11262) );
  NAND20 U74681 ( .A(N3400), .B(n65578), .Q(n66045) );
  CLKIN0 U74682 ( .A(n66045), .Q(\r37771/carry [4]) );
  NAND20 U74683 ( .A(N3364), .B(n65578), .Q(n66046) );
  CLKIN0 U74684 ( .A(n66046), .Q(\r40768/carry [4]) );
  NAND20 U74685 ( .A(N3382), .B(n65584), .Q(n66047) );
  CLKIN0 U74686 ( .A(n66047), .Q(\r32400/carry [4]) );
  NAND20 U74687 ( .A(N5515), .B(n65578), .Q(n66048) );
  CLKIN0 U74688 ( .A(n66048), .Q(\add_0_root_sub_0_root_sub_375_7/carry [4])
         );
  NAND20 U74689 ( .A(N3209), .B(n65584), .Q(n66049) );
  CLKIN0 U74690 ( .A(n66049), .Q(\r31798/carry [4]) );
  NAND20 U74691 ( .A(N3227), .B(n65578), .Q(n66050) );
  CLKIN0 U74692 ( .A(n66050), .Q(\r36567/carry [4]) );
  XNR20 U74693 ( .A(n65601), .B(\r12189/carry[5] ), .Q(N11290) );
  NOR20 U74694 ( .A(\r12189/carry[4] ), .B(n65599), .Q(n66051) );
  XNR20 U74695 ( .A(\r12189/carry[4] ), .B(n65598), .Q(N11291) );
  CLKIN0 U74696 ( .A(n66051), .Q(\r12189/carry[5] ) );
  NAND20 U74697 ( .A(N11292), .B(n65584), .Q(n66052) );
  CLKIN0 U74698 ( .A(n66052), .Q(\r12191/carry [4]) );
  NOR20 U74699 ( .A(\r12189/carry[3] ), .B(n65594), .Q(n66053) );
  XNR20 U74700 ( .A(\r12189/carry[3] ), .B(n65594), .Q(N11292) );
  CLKIN0 U74701 ( .A(n66053), .Q(\r12189/carry[4] ) );
  NOR20 U74702 ( .A(\add_1_root_add_0_root_sub_328_8_cf/carry[2] ), .B(N1167), 
        .Q(n66054) );
  CLKIN0 U74703 ( .A(n66054), .Q(\r12189/carry[3] ) );
  XNR20 U74704 ( .A(n65601), .B(\r12188/carry [5]), .Q(N11284) );
  NOR20 U74705 ( .A(\r12188/carry [4]), .B(n65599), .Q(n66055) );
  XNR20 U74706 ( .A(\r12188/carry [4]), .B(n65598), .Q(N11285) );
  CLKIN0 U74707 ( .A(n66055), .Q(\r12188/carry [5]) );
  NAND20 U74708 ( .A(N11286), .B(n65580), .Q(n66056) );
  CLKIN0 U74709 ( .A(n66056), .Q(\r12190/carry [4]) );
  NOR20 U74710 ( .A(\r34786/carry [3]), .B(n65594), .Q(n66057) );
  XNR20 U74711 ( .A(\r34786/carry [3]), .B(n65594), .Q(N11286) );
  NAND20 U74712 ( .A(N5206), .B(n65578), .Q(n66058) );
  CLKIN0 U74713 ( .A(n66058), .Q(\add_0_root_sub_0_root_sub_369_9/carry [4])
         );
  NAND20 U74714 ( .A(N5170), .B(n65578), .Q(n66059) );
  CLKIN0 U74715 ( .A(n66059), .Q(\add_0_root_sub_0_root_sub_369_3/carry [4])
         );
  NAND20 U74716 ( .A(N5188), .B(n65580), .Q(n66060) );
  CLKIN0 U74717 ( .A(n66060), .Q(\add_0_root_sub_0_root_sub_369_6/carry [4])
         );
  NAND20 U74718 ( .A(N5360), .B(n65584), .Q(n66061) );
  CLKIN0 U74719 ( .A(n66061), .Q(\add_0_root_sub_0_root_sub_372_8/carry [4])
         );
  NAND20 U74720 ( .A(N3054), .B(n65578), .Q(n66062) );
  CLKIN0 U74721 ( .A(n66062), .Q(\r37169/carry [4]) );
  NAND20 U74722 ( .A(N5342), .B(n65578), .Q(n66063) );
  CLKIN0 U74723 ( .A(n66063), .Q(\add_0_root_sub_0_root_sub_372_5/carry [4])
         );
  NOR20 U74724 ( .A(\sub_1_root_sub_0_root_sub_136_2/A[4] ), .B(n65420), .Q(
        n66065) );
  NOR20 U74725 ( .A(n66069), .B(N1367), .Q(n66064) );
  NOR20 U74726 ( .A(n66070), .B(N1368), .Q(n66067) );
  OAI210 U74727 ( .A(n65741), .B(n66857), .C(n66069), .Q(N1376) );
  OAI210 U74728 ( .A(n66065), .B(n66480), .C(n66070), .Q(N1377) );
  AOI210 U74729 ( .A(n66070), .B(N1368), .C(n66067), .Q(n66066) );
  NOR20 U74730 ( .A(N1371), .B(n66071), .Q(n66068) );
  CLKIN0 U74731 ( .A(n66072), .Q(n66071) );
  OAI210 U74732 ( .A(n66067), .B(n66073), .C(n66072), .Q(N1379) );
  NAND20 U74733 ( .A(n66072), .B(n66073), .Q(N1403) );
  NAND20 U74734 ( .A(n66067), .B(n66073), .Q(n66072) );
  CLKIN0 U74735 ( .A(N1371), .Q(n66073) );
  NOR20 U74736 ( .A(\sub_1_root_sub_0_root_sub_167_2/A[4] ), .B(n65511), .Q(
        n66075) );
  NOR20 U74737 ( .A(n66079), .B(N1910), .Q(n66074) );
  NOR20 U74738 ( .A(n66080), .B(N1911), .Q(n66077) );
  OAI210 U74739 ( .A(n65740), .B(n66871), .C(n66079), .Q(N1919) );
  OAI210 U74740 ( .A(n66075), .B(n66645), .C(n66080), .Q(N1920) );
  AOI210 U74741 ( .A(n66080), .B(N1911), .C(n66077), .Q(n66076) );
  NOR20 U74742 ( .A(N1914), .B(n66081), .Q(n66078) );
  CLKIN0 U74743 ( .A(n66082), .Q(n66081) );
  OAI210 U74744 ( .A(n66077), .B(n66083), .C(n66082), .Q(N1922) );
  NAND20 U74745 ( .A(n66077), .B(n66083), .Q(n66082) );
  CLKIN0 U74746 ( .A(N1914), .Q(n66083) );
  NOR20 U74747 ( .A(n66103), .B(N1167), .Q(n66085) );
  AOI210 U74748 ( .A(n66103), .B(n65916), .C(n66085), .Q(n66084) );
  NAND20 U74749 ( .A(n66085), .B(n65595), .Q(n66086) );
  OAI210 U74750 ( .A(n66085), .B(n65595), .C(n66086), .Q(N3364) );
  XNR20 U74751 ( .A(n65599), .B(n66086), .Q(N3365) );
  NOR20 U74752 ( .A(n66086), .B(n65599), .Q(n66087) );
  XOR20 U74753 ( .A(n66087), .B(n[5]), .Q(N3366) );
  NOR20 U74754 ( .A(n66103), .B(N1167), .Q(n66089) );
  AOI210 U74755 ( .A(n66097), .B(n65918), .C(n66089), .Q(n66088) );
  NAND20 U74756 ( .A(n66089), .B(n65596), .Q(n66090) );
  OAI210 U74757 ( .A(n66089), .B(n65595), .C(n66090), .Q(N3400) );
  XNR20 U74758 ( .A(n65599), .B(n66090), .Q(N3401) );
  NOR20 U74759 ( .A(n66090), .B(n65599), .Q(n66091) );
  XOR20 U74760 ( .A(n66091), .B(n[5]), .Q(N3402) );
  NOR20 U74761 ( .A(n65745), .B(n65889), .Q(n66092) );
  OAI210 U74762 ( .A(n65808), .B(n65771), .C(n66097), .Q(N998) );
  NOR20 U74763 ( .A(n66097), .B(N1167), .Q(n66094) );
  AOI210 U74764 ( .A(n66097), .B(n65917), .C(n66094), .Q(n66093) );
  NAND20 U74765 ( .A(n66094), .B(n65595), .Q(n66095) );
  OAI210 U74766 ( .A(n66094), .B(n65595), .C(n66095), .Q(N3054) );
  XNR20 U74767 ( .A(n65599), .B(n66095), .Q(N3055) );
  NOR20 U74768 ( .A(n66095), .B(n[4]), .Q(n66096) );
  XOR20 U74769 ( .A(n66096), .B(n65601), .Q(N3056) );
  NOR20 U74770 ( .A(n65755), .B(n65871), .Q(n66098) );
  OAI210 U74771 ( .A(n65791), .B(n65759), .C(n66103), .Q(N1022) );
  NOR20 U74772 ( .A(n66103), .B(N1167), .Q(n66100) );
  AOI210 U74773 ( .A(n66103), .B(n65916), .C(n66100), .Q(n66099) );
  NAND20 U74774 ( .A(n66100), .B(n65596), .Q(n66101) );
  OAI210 U74775 ( .A(n66100), .B(n65596), .C(n66101), .Q(N3227) );
  XNR20 U74776 ( .A(n65599), .B(n66101), .Q(N3228) );
  NOR20 U74777 ( .A(n66101), .B(n65599), .Q(n66102) );
  XOR20 U74778 ( .A(n66102), .B(n65601), .Q(N3229) );
  XOR20 U74779 ( .A(\r32997/carry [5]), .B(N11428), .Q(N1188) );
  NOR20 U74780 ( .A(N1208), .B(n65903), .Q(n66109) );
  NOR20 U74781 ( .A(n66114), .B(N1167), .Q(n66111) );
  AOI210 U74782 ( .A(n66114), .B(n65918), .C(n66111), .Q(n66110) );
  NAND20 U74783 ( .A(n66111), .B(n65595), .Q(n66112) );
  OAI210 U74784 ( .A(n66111), .B(n65596), .C(n66112), .Q(N3382) );
  XNR20 U74785 ( .A(n65599), .B(n66112), .Q(N3383) );
  NOR20 U74786 ( .A(n66112), .B(n[4]), .Q(n66113) );
  XOR20 U74787 ( .A(n66113), .B(n65601), .Q(N3384) );
  OAI210 U74788 ( .A(n65787), .B(n65761), .C(n66103), .Q(N1016) );
  NOR20 U74789 ( .A(n66097), .B(N1167), .Q(n66116) );
  AOI210 U74790 ( .A(n66114), .B(n65916), .C(n66116), .Q(n66115) );
  NAND20 U74791 ( .A(n66116), .B(n65596), .Q(n66117) );
  OAI210 U74792 ( .A(n66116), .B(n65595), .C(n66117), .Q(N3209) );
  XNR20 U74793 ( .A(n65599), .B(n66117), .Q(N3210) );
  NOR20 U74794 ( .A(n66117), .B(n[4]), .Q(n66118) );
  XOR20 U74795 ( .A(n66118), .B(n65601), .Q(N3211) );
  XOR20 U74796 ( .A(\r31196/carry [5]), .B(N11410), .Q(N1176) );
  XOR20 U74797 ( .A(\sub_420_6_cf/carry [5]), .B(N11524), .Q(N1260) );
  XOR20 U74798 ( .A(\sub_348_6_cf/carry [5]), .B(N11536), .Q(N972) );
  XOR20 U74799 ( .A(\sub_417_9_cf/carry [5]), .B(N11506), .Q(N1248) );
  XOR20 U74800 ( .A(\sub_345_9_cf/carry [5]), .B(N11518), .Q(N960) );
  XOR20 U74801 ( .A(\r13451/carry [5]), .B(N1122), .Q(N1116) );
  NOR20 U74802 ( .A(n66097), .B(n65918), .Q(n66128) );
  AOI210 U74803 ( .A(n66103), .B(n65915), .C(n66128), .Q(n66127) );
  NAND20 U74804 ( .A(n66128), .B(n65595), .Q(n66129) );
  OAI210 U74805 ( .A(n66128), .B(n65595), .C(n66129), .Q(N5515) );
  XNR20 U74806 ( .A(n65599), .B(n66129), .Q(N5516) );
  NOR20 U74807 ( .A(n66129), .B(n[4]), .Q(n66130) );
  XOR20 U74808 ( .A(n66130), .B(n[5]), .Q(N5517) );
  NOR20 U74809 ( .A(n66114), .B(N1167), .Q(n66132) );
  AOI210 U74810 ( .A(n66114), .B(N1167), .C(n66132), .Q(n66131) );
  NAND20 U74811 ( .A(n66132), .B(n65596), .Q(n66133) );
  OAI210 U74812 ( .A(n66132), .B(n65596), .C(n66133), .Q(N3245) );
  XNR20 U74813 ( .A(n65599), .B(n66133), .Q(N3246) );
  NOR20 U74814 ( .A(n66133), .B(n[4]), .Q(n66134) );
  XOR20 U74815 ( .A(n66134), .B(n[5]), .Q(N3247) );
  NOR20 U74816 ( .A(n66114), .B(n65918), .Q(n66136) );
  AOI210 U74817 ( .A(n66103), .B(n65917), .C(n66136), .Q(n66135) );
  NAND20 U74818 ( .A(n66136), .B(n65595), .Q(n66137) );
  OAI210 U74819 ( .A(n66136), .B(n65596), .C(n66137), .Q(N5360) );
  XNR20 U74820 ( .A(n65599), .B(n66137), .Q(N5361) );
  NOR20 U74821 ( .A(n66137), .B(n[4]), .Q(n66138) );
  XOR20 U74822 ( .A(n66138), .B(n[5]), .Q(N5362) );
  NOR20 U74823 ( .A(n66103), .B(n65917), .Q(n66140) );
  AOI210 U74824 ( .A(n66103), .B(n65918), .C(n66140), .Q(n66139) );
  NAND20 U74825 ( .A(n66140), .B(n65596), .Q(n66141) );
  OAI210 U74826 ( .A(n66140), .B(n65595), .C(n66141), .Q(N5342) );
  XNR20 U74827 ( .A(n65599), .B(n66141), .Q(N5343) );
  NOR20 U74828 ( .A(n66141), .B(n[4]), .Q(n66142) );
  XOR20 U74829 ( .A(n66142), .B(n[5]), .Q(N5344) );
  NOR20 U74830 ( .A(n66103), .B(n65916), .Q(n66144) );
  AOI210 U74831 ( .A(n66097), .B(N1167), .C(n66144), .Q(n66143) );
  NAND20 U74832 ( .A(n66144), .B(n65595), .Q(n66145) );
  OAI210 U74833 ( .A(n66144), .B(n65595), .C(n66145), .Q(N3090) );
  XNR20 U74834 ( .A(n65599), .B(n66145), .Q(N3091) );
  NOR20 U74835 ( .A(n66145), .B(n[4]), .Q(n66146) );
  XOR20 U74836 ( .A(n66146), .B(n65601), .Q(N3092) );
  NOR20 U74837 ( .A(n66097), .B(N1167), .Q(n66148) );
  AOI210 U74838 ( .A(n66103), .B(n65918), .C(n66148), .Q(n66147) );
  NAND20 U74839 ( .A(n66148), .B(n65595), .Q(n66149) );
  OAI210 U74840 ( .A(n66148), .B(n65596), .C(n66149), .Q(N3072) );
  XNR20 U74841 ( .A(n65599), .B(n66149), .Q(N3073) );
  NOR20 U74842 ( .A(n66149), .B(n[4]), .Q(n66150) );
  XOR20 U74843 ( .A(n66150), .B(n65601), .Q(N3074) );
  NOR20 U74844 ( .A(n66114), .B(N1167), .Q(n66152) );
  AOI210 U74845 ( .A(n66114), .B(n65915), .C(n66152), .Q(n66151) );
  NAND20 U74846 ( .A(n66152), .B(n65596), .Q(n66153) );
  OAI210 U74847 ( .A(n66152), .B(n65596), .C(n66153), .Q(N5206) );
  XNR20 U74848 ( .A(n65599), .B(n66153), .Q(N5207) );
  NOR20 U74849 ( .A(n66153), .B(n[4]), .Q(n66154) );
  XOR20 U74850 ( .A(n66154), .B(n[5]), .Q(N5208) );
  NOR20 U74851 ( .A(n66097), .B(N1167), .Q(n66156) );
  AOI210 U74852 ( .A(n66103), .B(n65917), .C(n66156), .Q(n66155) );
  NAND20 U74853 ( .A(n66156), .B(n65595), .Q(n66157) );
  OAI210 U74854 ( .A(n66156), .B(n65596), .C(n66157), .Q(N5188) );
  XNR20 U74855 ( .A(n65599), .B(n66157), .Q(N5189) );
  NOR20 U74856 ( .A(n66157), .B(n[4]), .Q(n66158) );
  XOR20 U74857 ( .A(n66158), .B(n65601), .Q(N5190) );
  NOR20 U74858 ( .A(n66114), .B(N1167), .Q(n66160) );
  AOI210 U74859 ( .A(n66114), .B(N1167), .C(n66160), .Q(n66159) );
  NAND20 U74860 ( .A(n66160), .B(n65596), .Q(n66161) );
  OAI210 U74861 ( .A(n66160), .B(n65595), .C(n66161), .Q(N5170) );
  XNR20 U74862 ( .A(n65599), .B(n66161), .Q(N5171) );
  NOR20 U74863 ( .A(n66161), .B(n[4]), .Q(n66162) );
  XOR20 U74864 ( .A(n66162), .B(n65601), .Q(N5172) );
  NOR20 U74865 ( .A(n66097), .B(N1167), .Q(n66164) );
  AOI210 U74866 ( .A(n66097), .B(n65915), .C(n66164), .Q(n66163) );
  NAND20 U74867 ( .A(n66164), .B(n65596), .Q(n66165) );
  OAI210 U74868 ( .A(n66164), .B(n65596), .C(n66165), .Q(N2936) );
  XNR20 U74869 ( .A(n65599), .B(n66165), .Q(N2937) );
  NOR20 U74870 ( .A(n66165), .B(n[4]), .Q(n66166) );
  XOR20 U74871 ( .A(n66166), .B(n[5]), .Q(N2938) );
  XNR20 U74872 ( .A(N2913), .B(n65581), .Q(N2919) );
  NAND20 U74873 ( .A(n65579), .B(N2919), .Q(n66167) );
  IMUX20 U74874 ( .A(n66167), .B(n66168), .S(N2914), .Q(N2920) );
  XNR20 U74875 ( .A(n65605), .B(n65578), .Q(N2901) );
  NAND20 U74876 ( .A(n65584), .B(N2901), .Q(n66169) );
  IMUX20 U74877 ( .A(n66169), .B(n66170), .S(N2896), .Q(N2902) );
  XNR22 U74878 ( .A(n65602), .B(n65578), .Q(N3510) );
  XNR22 U74879 ( .A(n65602), .B(n65578), .Q(N3637) );
  OAI212 U74880 ( .A(n66717), .B(n66716), .C(n66643), .Q(N3760) );
  OAI212 U74881 ( .A(n66727), .B(n66726), .C(n66643), .Q(N4021) );
  OAI212 U74882 ( .A(n66760), .B(n66759), .C(n66643), .Q(N4297) );
  OAI212 U74883 ( .A(n66782), .B(n66781), .C(n66643), .Q(N4436) );
  OAI212 U74884 ( .A(n66792), .B(n66791), .C(n66643), .Q(N4573) );
  OAI212 U74885 ( .A(n66823), .B(n66822), .C(n66643), .Q(N4849) );
  OAI212 U74886 ( .A(n66845), .B(n66844), .C(n66643), .Q(N4988) );
  OAI212 U74887 ( .A(n66856), .B(n66855), .C(n66643), .Q(N5124) );
  OAI212 U74888 ( .A(n66858), .B(n66481), .C(n66859), .Q(N1367) );
  OAI212 U74889 ( .A(n65546), .B(N1301), .C(N1302), .Q(n66867) );
  OAI212 U74890 ( .A(n66870), .B(n66869), .C(n66482), .Q(N1560) );
  OAI212 U74891 ( .A(n66872), .B(n66646), .C(n66873), .Q(N1910) );
  OAI212 U74892 ( .A(N1843), .B(N1844), .C(N1845), .Q(n66881) );
  OAI212 U74893 ( .A(n66884), .B(n66883), .C(n66570), .Q(N2103) );
  OAI222 U74894 ( .A(N1294), .B(N1295), .C(n66540), .D(N1295), .Q(N1503) );
  OAI222 U74895 ( .A(N1837), .B(N1838), .C(n66647), .D(N1838), .Q(N2046) );
endmodule


module Connect4_DW01_add_96 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [31:1] carry;

  ADD32 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADD32 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADD32 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADD32 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADD32 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADD32 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADD32 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADD32 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADD32 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADD32 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADD32 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADD32 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADD32 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADD32 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADD32 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADD32 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADD32 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADD32 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADD32 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADD32 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADD32 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADD32 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADD32 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR31 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Q(SUM[31]) );
  INV3 U1 ( .A(n2), .Q(carry[3]) );
  NOR21 U2 ( .A(B[2]), .B(carry[2]), .Q(n2) );
  INV3 U3 ( .A(B[0]), .Q(SUM[0]) );
  INV3 U4 ( .A(n1), .Q(carry[2]) );
  NOR21 U5 ( .A(B[1]), .B(B[0]), .Q(n1) );
  XNR22 U6 ( .A(B[0]), .B(B[1]), .Q(SUM[1]) );
  XNR22 U7 ( .A(carry[2]), .B(B[2]), .Q(SUM[2]) );
endmodule


module Connect4_DW01_add_97 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [31:1] carry;

  ADD32 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADD32 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADD32 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADD32 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADD32 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADD32 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADD32 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADD32 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADD32 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADD32 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADD32 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADD32 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADD32 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADD32 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADD32 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADD32 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADD32 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADD32 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADD32 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADD32 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADD32 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADD32 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADD32 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR31 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Q(SUM[31]) );
  INV3 U1 ( .A(n2), .Q(carry[3]) );
  NOR21 U2 ( .A(B[2]), .B(carry[2]), .Q(n2) );
  INV3 U3 ( .A(B[0]), .Q(SUM[0]) );
  INV3 U4 ( .A(n1), .Q(carry[2]) );
  NOR21 U5 ( .A(B[1]), .B(B[0]), .Q(n1) );
  XNR22 U6 ( .A(B[0]), .B(B[1]), .Q(SUM[1]) );
  XNR22 U7 ( .A(carry[2]), .B(B[2]), .Q(SUM[2]) );
endmodule

